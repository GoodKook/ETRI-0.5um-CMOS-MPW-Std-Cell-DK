magic
tech scmos
magscale 1 2
timestamp 1746272870
<< nwell >>
rect 2409 4436 2445 4440
rect -2 4224 4782 4436
rect -2 3744 4782 3956
rect 2009 3740 2045 3744
rect 3669 3476 3705 3480
rect -2 3382 4782 3476
rect -3 3264 4783 3382
rect 1515 3260 1551 3264
rect -2 2784 4782 2996
rect 2829 2516 2865 2520
rect -2 2304 4782 2516
rect 3669 2300 3705 2304
rect 2589 2036 2625 2040
rect -2 1918 4783 2036
rect -2 1824 4782 1918
rect 4109 1820 4145 1824
rect -2 1344 4782 1556
rect 2329 1340 2365 1344
rect -2 864 4782 1076
rect -2 502 4782 596
rect -2 384 4783 502
rect 3589 380 3625 384
rect -2 -2 4782 116
<< ntransistor >>
rect 52 4536 56 4556
rect 74 4516 78 4556
rect 82 4516 86 4556
rect 168 4496 172 4556
rect 176 4496 180 4556
rect 184 4496 188 4556
rect 232 4496 236 4556
rect 240 4496 244 4556
rect 248 4496 252 4556
rect 368 4496 372 4556
rect 376 4496 380 4556
rect 384 4496 388 4556
rect 434 4516 438 4556
rect 442 4516 446 4556
rect 464 4536 468 4556
rect 531 4516 535 4556
rect 551 4516 555 4556
rect 571 4516 575 4556
rect 631 4516 635 4556
rect 651 4516 655 4556
rect 671 4516 675 4556
rect 768 4496 772 4556
rect 776 4496 780 4556
rect 784 4496 788 4556
rect 832 4496 836 4556
rect 840 4496 844 4556
rect 848 4496 852 4556
rect 933 4516 937 4556
rect 943 4516 947 4556
rect 1012 4496 1016 4556
rect 1020 4496 1024 4556
rect 1028 4496 1032 4556
rect 1114 4516 1118 4556
rect 1122 4516 1126 4556
rect 1144 4536 1148 4556
rect 1233 4516 1237 4556
rect 1243 4516 1247 4556
rect 1305 4536 1309 4556
rect 1325 4536 1329 4556
rect 1385 4516 1389 4556
rect 1405 4516 1409 4556
rect 1425 4516 1429 4556
rect 1493 4516 1497 4556
rect 1503 4516 1507 4556
rect 1551 4536 1555 4556
rect 1571 4536 1575 4556
rect 1632 4496 1636 4556
rect 1640 4496 1644 4556
rect 1648 4496 1652 4556
rect 1752 4536 1756 4556
rect 1774 4516 1778 4556
rect 1782 4516 1786 4556
rect 1831 4536 1835 4556
rect 1905 4536 1909 4556
rect 1954 4516 1958 4556
rect 1962 4516 1966 4556
rect 1984 4536 1988 4556
rect 2051 4536 2055 4556
rect 2071 4536 2075 4556
rect 2131 4536 2135 4556
rect 2191 4516 2195 4556
rect 2211 4516 2215 4556
rect 2231 4516 2235 4556
rect 2305 4516 2309 4556
rect 2325 4516 2329 4556
rect 2345 4516 2349 4556
rect 2365 4516 2369 4556
rect 2411 4536 2415 4556
rect 2431 4536 2435 4556
rect 2451 4516 2455 4556
rect 2514 4516 2518 4556
rect 2522 4516 2526 4556
rect 2544 4536 2548 4556
rect 2646 4516 2650 4556
rect 2654 4516 2658 4556
rect 2674 4516 2678 4556
rect 2682 4516 2686 4556
rect 2735 4516 2739 4556
rect 2755 4536 2759 4556
rect 2765 4536 2769 4556
rect 2787 4536 2791 4556
rect 2797 4536 2801 4556
rect 2819 4536 2823 4556
rect 2865 4536 2869 4556
rect 2873 4536 2877 4556
rect 2893 4536 2897 4556
rect 2903 4536 2907 4556
rect 2925 4516 2929 4556
rect 2985 4536 2989 4556
rect 3045 4516 3049 4556
rect 3065 4516 3069 4556
rect 3085 4516 3089 4556
rect 3145 4536 3149 4556
rect 3165 4536 3169 4556
rect 3225 4516 3229 4556
rect 3245 4516 3249 4556
rect 3265 4516 3269 4556
rect 3325 4536 3329 4556
rect 3345 4536 3349 4556
rect 3405 4536 3409 4556
rect 3451 4516 3455 4556
rect 3473 4536 3477 4556
rect 3483 4536 3487 4556
rect 3503 4536 3507 4556
rect 3511 4536 3515 4556
rect 3557 4536 3561 4556
rect 3579 4536 3583 4556
rect 3589 4536 3593 4556
rect 3611 4536 3615 4556
rect 3621 4536 3625 4556
rect 3641 4516 3645 4556
rect 3691 4516 3695 4556
rect 3711 4516 3715 4556
rect 3731 4516 3735 4556
rect 3793 4516 3797 4556
rect 3803 4516 3807 4556
rect 3885 4516 3889 4556
rect 3905 4516 3909 4556
rect 3925 4516 3929 4556
rect 3945 4516 3949 4556
rect 3965 4516 3969 4556
rect 3985 4516 3989 4556
rect 4005 4516 4009 4556
rect 4025 4516 4029 4556
rect 4083 4516 4087 4556
rect 4105 4536 4109 4556
rect 4153 4516 4157 4556
rect 4163 4516 4167 4556
rect 4231 4536 4235 4556
rect 4291 4516 4295 4556
rect 4311 4516 4315 4556
rect 4331 4516 4335 4556
rect 4391 4516 4395 4556
rect 4413 4536 4417 4556
rect 4423 4536 4427 4556
rect 4443 4536 4447 4556
rect 4451 4536 4455 4556
rect 4497 4536 4501 4556
rect 4519 4536 4523 4556
rect 4529 4536 4533 4556
rect 4551 4536 4555 4556
rect 4561 4536 4565 4556
rect 4581 4516 4585 4556
rect 4631 4536 4635 4556
rect 4653 4516 4657 4556
rect 4713 4516 4717 4556
rect 4723 4516 4727 4556
rect 53 4104 57 4144
rect 63 4104 67 4144
rect 114 4104 118 4144
rect 122 4104 126 4144
rect 144 4104 148 4124
rect 233 4104 237 4144
rect 243 4104 247 4144
rect 305 4104 309 4124
rect 325 4104 329 4124
rect 385 4104 389 4144
rect 405 4104 409 4144
rect 425 4104 429 4144
rect 471 4104 475 4144
rect 491 4104 495 4144
rect 511 4104 515 4144
rect 585 4104 589 4124
rect 652 4104 656 4124
rect 674 4104 678 4144
rect 682 4104 686 4144
rect 745 4104 749 4124
rect 792 4104 796 4164
rect 800 4104 804 4164
rect 808 4104 812 4164
rect 926 4104 930 4144
rect 934 4104 938 4144
rect 954 4104 958 4144
rect 962 4104 966 4144
rect 1048 4104 1052 4164
rect 1056 4104 1060 4164
rect 1064 4104 1068 4164
rect 1112 4104 1116 4164
rect 1120 4104 1124 4164
rect 1128 4104 1132 4164
rect 1233 4104 1237 4144
rect 1243 4104 1247 4144
rect 1328 4104 1332 4164
rect 1336 4104 1340 4164
rect 1344 4104 1348 4164
rect 1413 4104 1417 4144
rect 1423 4104 1427 4144
rect 1472 4104 1476 4164
rect 1480 4104 1484 4164
rect 1488 4104 1492 4164
rect 1585 4104 1589 4124
rect 1605 4104 1609 4124
rect 1665 4104 1669 4124
rect 1685 4104 1689 4124
rect 1731 4104 1735 4144
rect 1751 4104 1755 4144
rect 1771 4104 1775 4144
rect 1853 4104 1857 4144
rect 1863 4104 1867 4144
rect 1911 4104 1915 4124
rect 1972 4104 1976 4164
rect 1980 4104 1984 4164
rect 1988 4104 1992 4164
rect 2072 4104 2076 4164
rect 2080 4104 2084 4164
rect 2088 4104 2092 4164
rect 2175 4104 2179 4144
rect 2195 4104 2199 4124
rect 2205 4104 2209 4124
rect 2227 4104 2231 4124
rect 2237 4104 2241 4124
rect 2259 4104 2263 4124
rect 2305 4104 2309 4124
rect 2313 4104 2317 4124
rect 2333 4104 2337 4124
rect 2343 4104 2347 4124
rect 2365 4104 2369 4144
rect 2411 4104 2415 4124
rect 2433 4104 2437 4144
rect 2505 4104 2509 4124
rect 2565 4104 2569 4124
rect 2585 4104 2589 4124
rect 2631 4104 2635 4144
rect 2653 4104 2657 4124
rect 2663 4104 2667 4124
rect 2683 4104 2687 4124
rect 2691 4104 2695 4124
rect 2737 4104 2741 4124
rect 2759 4104 2763 4124
rect 2769 4104 2773 4124
rect 2791 4104 2795 4124
rect 2801 4104 2805 4124
rect 2821 4104 2825 4144
rect 2871 4104 2875 4124
rect 2945 4104 2949 4124
rect 2965 4104 2969 4124
rect 3011 4104 3015 4144
rect 3031 4104 3035 4144
rect 3051 4104 3055 4144
rect 3113 4104 3117 4144
rect 3123 4104 3127 4144
rect 3213 4104 3217 4144
rect 3223 4104 3227 4144
rect 3293 4104 3297 4144
rect 3303 4104 3307 4144
rect 3351 4104 3355 4124
rect 3371 4104 3375 4124
rect 3435 4104 3439 4144
rect 3455 4104 3459 4124
rect 3465 4104 3469 4124
rect 3487 4104 3491 4124
rect 3497 4104 3501 4124
rect 3519 4104 3523 4124
rect 3565 4104 3569 4124
rect 3573 4104 3577 4124
rect 3593 4104 3597 4124
rect 3603 4104 3607 4124
rect 3625 4104 3629 4144
rect 3693 4104 3697 4144
rect 3703 4104 3707 4144
rect 3751 4104 3755 4124
rect 3771 4104 3775 4124
rect 3831 4104 3835 4144
rect 3853 4104 3857 4124
rect 3863 4104 3867 4124
rect 3883 4104 3887 4124
rect 3891 4104 3895 4124
rect 3937 4104 3941 4124
rect 3959 4104 3963 4124
rect 3969 4104 3973 4124
rect 3991 4104 3995 4124
rect 4001 4104 4005 4124
rect 4021 4104 4025 4144
rect 4071 4104 4075 4124
rect 4091 4104 4095 4124
rect 4172 4104 4176 4124
rect 4194 4104 4198 4144
rect 4202 4104 4206 4144
rect 4251 4104 4255 4124
rect 4273 4104 4277 4144
rect 4345 4104 4349 4124
rect 4365 4104 4369 4124
rect 4432 4104 4436 4124
rect 4454 4104 4458 4144
rect 4462 4104 4466 4144
rect 4511 4104 4515 4144
rect 4533 4104 4537 4124
rect 4543 4104 4547 4124
rect 4563 4104 4567 4124
rect 4571 4104 4575 4124
rect 4617 4104 4621 4124
rect 4639 4104 4643 4124
rect 4649 4104 4653 4124
rect 4671 4104 4675 4124
rect 4681 4104 4685 4124
rect 4701 4104 4705 4144
rect 53 4036 57 4076
rect 63 4036 67 4076
rect 113 4036 117 4076
rect 123 4036 127 4076
rect 213 4036 217 4076
rect 223 4036 227 4076
rect 285 4036 289 4076
rect 305 4036 309 4076
rect 325 4036 329 4076
rect 374 4036 378 4076
rect 382 4036 386 4076
rect 404 4056 408 4076
rect 485 4056 489 4076
rect 505 4056 509 4076
rect 553 4036 557 4076
rect 563 4036 567 4076
rect 631 4036 635 4076
rect 651 4036 655 4076
rect 671 4036 675 4076
rect 768 4016 772 4076
rect 776 4016 780 4076
rect 784 4016 788 4076
rect 832 4016 836 4076
rect 840 4016 844 4076
rect 848 4016 852 4076
rect 945 4036 949 4076
rect 965 4036 969 4076
rect 985 4036 989 4076
rect 1031 4036 1035 4076
rect 1051 4036 1055 4076
rect 1071 4036 1075 4076
rect 1145 4056 1149 4076
rect 1228 4016 1232 4076
rect 1236 4016 1240 4076
rect 1244 4016 1248 4076
rect 1291 4056 1295 4076
rect 1352 4016 1356 4076
rect 1360 4016 1364 4076
rect 1368 4016 1372 4076
rect 1452 4016 1456 4076
rect 1460 4016 1464 4076
rect 1468 4016 1472 4076
rect 1553 4036 1557 4076
rect 1563 4036 1567 4076
rect 1645 4056 1649 4076
rect 1665 4056 1669 4076
rect 1735 4036 1739 4076
rect 1755 4036 1759 4076
rect 1765 4036 1769 4076
rect 1825 4036 1829 4076
rect 1845 4036 1849 4076
rect 1865 4036 1869 4076
rect 1911 4056 1915 4076
rect 1931 4056 1935 4076
rect 2005 4056 2009 4076
rect 2051 4036 2055 4076
rect 2071 4036 2075 4076
rect 2091 4036 2095 4076
rect 2151 4056 2155 4076
rect 2213 4036 2217 4076
rect 2223 4036 2227 4076
rect 2292 4016 2296 4076
rect 2300 4016 2304 4076
rect 2308 4016 2312 4076
rect 2391 4056 2395 4076
rect 2413 4036 2417 4076
rect 2471 4036 2475 4076
rect 2491 4036 2495 4076
rect 2511 4036 2515 4076
rect 2531 4036 2535 4076
rect 2551 4036 2555 4076
rect 2571 4036 2575 4076
rect 2591 4036 2595 4076
rect 2611 4036 2615 4076
rect 2675 4036 2679 4076
rect 2695 4056 2699 4076
rect 2705 4056 2709 4076
rect 2727 4056 2731 4076
rect 2737 4056 2741 4076
rect 2759 4056 2763 4076
rect 2805 4056 2809 4076
rect 2813 4056 2817 4076
rect 2833 4056 2837 4076
rect 2843 4056 2847 4076
rect 2865 4036 2869 4076
rect 2911 4056 2915 4076
rect 2971 4036 2975 4076
rect 2991 4036 2995 4076
rect 3011 4036 3015 4076
rect 3071 4056 3075 4076
rect 3091 4056 3095 4076
rect 3153 4036 3157 4076
rect 3163 4036 3167 4076
rect 3252 4056 3256 4076
rect 3274 4036 3278 4076
rect 3282 4036 3286 4076
rect 3331 4036 3335 4076
rect 3341 4036 3345 4076
rect 3361 4036 3365 4076
rect 3445 4056 3449 4076
rect 3465 4056 3469 4076
rect 3525 4056 3529 4076
rect 3571 4036 3575 4076
rect 3593 4056 3597 4076
rect 3603 4056 3607 4076
rect 3623 4056 3627 4076
rect 3631 4056 3635 4076
rect 3677 4056 3681 4076
rect 3699 4056 3703 4076
rect 3709 4056 3713 4076
rect 3731 4056 3735 4076
rect 3741 4056 3745 4076
rect 3761 4036 3765 4076
rect 3832 4056 3836 4076
rect 3854 4036 3858 4076
rect 3862 4036 3866 4076
rect 3911 4056 3915 4076
rect 3931 4056 3935 4076
rect 4005 4056 4009 4076
rect 4025 4056 4029 4076
rect 4071 4036 4075 4076
rect 4081 4036 4085 4076
rect 4101 4036 4105 4076
rect 4171 4036 4175 4076
rect 4191 4036 4195 4076
rect 4211 4036 4215 4076
rect 4285 4036 4289 4076
rect 4305 4036 4309 4076
rect 4325 4036 4329 4076
rect 4385 4056 4389 4076
rect 4431 4036 4435 4076
rect 4453 4056 4457 4076
rect 4463 4056 4467 4076
rect 4483 4056 4487 4076
rect 4491 4056 4495 4076
rect 4537 4056 4541 4076
rect 4559 4056 4563 4076
rect 4569 4056 4573 4076
rect 4591 4056 4595 4076
rect 4601 4056 4605 4076
rect 4621 4036 4625 4076
rect 4671 4056 4675 4076
rect 45 3624 49 3644
rect 65 3624 69 3644
rect 111 3624 115 3664
rect 131 3624 135 3664
rect 151 3624 155 3664
rect 225 3624 229 3644
rect 292 3624 296 3644
rect 314 3624 318 3664
rect 322 3624 326 3664
rect 395 3624 399 3664
rect 415 3624 419 3664
rect 425 3624 429 3664
rect 493 3624 497 3664
rect 503 3624 507 3664
rect 573 3624 577 3664
rect 583 3624 587 3664
rect 631 3624 635 3644
rect 691 3624 695 3664
rect 711 3624 715 3664
rect 731 3624 735 3664
rect 793 3624 797 3664
rect 803 3624 807 3664
rect 908 3624 912 3684
rect 916 3624 920 3684
rect 924 3624 928 3684
rect 974 3624 978 3664
rect 982 3624 986 3664
rect 1004 3624 1008 3644
rect 1072 3624 1076 3684
rect 1080 3624 1084 3684
rect 1088 3624 1092 3684
rect 1174 3624 1178 3664
rect 1182 3624 1186 3664
rect 1204 3624 1208 3644
rect 1271 3624 1275 3644
rect 1368 3624 1372 3684
rect 1376 3624 1380 3684
rect 1384 3624 1388 3684
rect 1445 3624 1449 3644
rect 1505 3624 1509 3664
rect 1525 3624 1529 3664
rect 1545 3624 1549 3664
rect 1605 3624 1609 3644
rect 1654 3624 1658 3664
rect 1662 3624 1666 3664
rect 1684 3624 1688 3644
rect 1751 3624 1755 3644
rect 1771 3624 1775 3644
rect 1852 3624 1856 3644
rect 1874 3624 1878 3664
rect 1882 3624 1886 3664
rect 1953 3624 1957 3664
rect 1963 3624 1967 3664
rect 2011 3624 2015 3644
rect 2031 3624 2035 3644
rect 2051 3624 2055 3664
rect 2111 3624 2115 3644
rect 2133 3624 2137 3664
rect 2205 3624 2209 3664
rect 2225 3624 2229 3664
rect 2245 3624 2249 3664
rect 2265 3624 2269 3664
rect 2285 3624 2289 3664
rect 2305 3624 2309 3664
rect 2325 3624 2329 3664
rect 2345 3624 2349 3664
rect 2395 3624 2399 3664
rect 2415 3624 2419 3644
rect 2425 3624 2429 3644
rect 2447 3624 2451 3644
rect 2457 3624 2461 3644
rect 2479 3624 2483 3644
rect 2525 3624 2529 3644
rect 2533 3624 2537 3644
rect 2553 3624 2557 3644
rect 2563 3624 2567 3644
rect 2585 3624 2589 3664
rect 2645 3624 2649 3664
rect 2665 3624 2669 3664
rect 2685 3624 2689 3664
rect 2745 3624 2749 3644
rect 2805 3624 2809 3644
rect 2825 3624 2829 3644
rect 2885 3624 2889 3644
rect 2905 3624 2909 3644
rect 2965 3624 2969 3644
rect 2985 3624 2989 3644
rect 3031 3624 3035 3644
rect 3105 3624 3109 3644
rect 3151 3624 3155 3664
rect 3171 3624 3175 3664
rect 3191 3624 3195 3664
rect 3272 3624 3276 3644
rect 3294 3624 3298 3664
rect 3302 3624 3306 3664
rect 3354 3624 3358 3664
rect 3362 3624 3366 3664
rect 3384 3624 3388 3644
rect 3451 3624 3455 3644
rect 3511 3624 3515 3664
rect 3521 3624 3525 3664
rect 3541 3624 3545 3664
rect 3611 3624 3615 3664
rect 3631 3624 3635 3664
rect 3651 3624 3655 3664
rect 3711 3624 3715 3664
rect 3731 3624 3735 3664
rect 3751 3624 3755 3664
rect 3815 3624 3819 3664
rect 3835 3624 3839 3644
rect 3845 3624 3849 3644
rect 3867 3624 3871 3644
rect 3877 3624 3881 3644
rect 3899 3624 3903 3644
rect 3945 3624 3949 3644
rect 3953 3624 3957 3644
rect 3973 3624 3977 3644
rect 3983 3624 3987 3644
rect 4005 3624 4009 3664
rect 4051 3624 4055 3644
rect 4073 3624 4077 3664
rect 4145 3624 4149 3644
rect 4165 3624 4169 3644
rect 4214 3624 4218 3664
rect 4222 3624 4226 3664
rect 4244 3624 4248 3644
rect 4311 3624 4315 3664
rect 4333 3624 4337 3644
rect 4343 3624 4347 3644
rect 4363 3624 4367 3644
rect 4371 3624 4375 3644
rect 4417 3624 4421 3644
rect 4439 3624 4443 3644
rect 4449 3624 4453 3644
rect 4471 3624 4475 3644
rect 4481 3624 4485 3644
rect 4501 3624 4505 3664
rect 4551 3624 4555 3644
rect 4573 3624 4577 3664
rect 4645 3624 4649 3644
rect 4691 3624 4695 3644
rect 53 3556 57 3596
rect 63 3556 67 3596
rect 115 3556 119 3596
rect 135 3576 139 3596
rect 145 3576 149 3596
rect 167 3576 171 3596
rect 177 3576 181 3596
rect 199 3576 203 3596
rect 245 3576 249 3596
rect 253 3576 257 3596
rect 273 3576 277 3596
rect 283 3576 287 3596
rect 305 3556 309 3596
rect 365 3576 369 3596
rect 433 3556 437 3596
rect 443 3556 447 3596
rect 505 3556 509 3596
rect 525 3556 529 3596
rect 545 3556 549 3596
rect 605 3556 609 3596
rect 625 3556 629 3596
rect 645 3556 649 3596
rect 693 3556 697 3596
rect 703 3556 707 3596
rect 771 3556 775 3596
rect 791 3556 795 3596
rect 811 3556 815 3596
rect 831 3556 835 3596
rect 891 3576 895 3596
rect 988 3536 992 3596
rect 996 3536 1000 3596
rect 1004 3536 1008 3596
rect 1054 3556 1058 3596
rect 1062 3556 1066 3596
rect 1084 3576 1088 3596
rect 1151 3576 1155 3596
rect 1171 3576 1175 3596
rect 1233 3556 1237 3596
rect 1243 3556 1247 3596
rect 1313 3556 1317 3596
rect 1323 3556 1327 3596
rect 1391 3556 1395 3596
rect 1411 3556 1415 3596
rect 1431 3556 1435 3596
rect 1495 3556 1499 3596
rect 1515 3576 1519 3596
rect 1525 3576 1529 3596
rect 1547 3576 1551 3596
rect 1557 3576 1561 3596
rect 1579 3576 1583 3596
rect 1625 3576 1629 3596
rect 1633 3576 1637 3596
rect 1653 3576 1657 3596
rect 1663 3576 1667 3596
rect 1685 3556 1689 3596
rect 1753 3556 1757 3596
rect 1763 3556 1767 3596
rect 1811 3556 1815 3596
rect 1831 3556 1835 3596
rect 1851 3556 1855 3596
rect 1911 3556 1915 3596
rect 1993 3556 1997 3596
rect 2003 3556 2007 3596
rect 2075 3556 2079 3596
rect 2095 3556 2099 3596
rect 2105 3556 2109 3596
rect 2153 3556 2157 3596
rect 2163 3556 2167 3596
rect 2232 3536 2236 3596
rect 2240 3536 2244 3596
rect 2248 3536 2252 3596
rect 2331 3576 2335 3596
rect 2391 3576 2395 3596
rect 2451 3556 2455 3596
rect 2473 3576 2477 3596
rect 2483 3576 2487 3596
rect 2503 3576 2507 3596
rect 2511 3576 2515 3596
rect 2557 3576 2561 3596
rect 2579 3576 2583 3596
rect 2589 3576 2593 3596
rect 2611 3576 2615 3596
rect 2621 3576 2625 3596
rect 2641 3556 2645 3596
rect 2691 3556 2695 3596
rect 2711 3556 2715 3596
rect 2731 3556 2735 3596
rect 2791 3576 2795 3596
rect 2813 3556 2817 3596
rect 2873 3556 2877 3596
rect 2883 3556 2887 3596
rect 2951 3556 2955 3596
rect 2973 3576 2977 3596
rect 2983 3576 2987 3596
rect 3003 3576 3007 3596
rect 3011 3576 3015 3596
rect 3057 3576 3061 3596
rect 3079 3576 3083 3596
rect 3089 3576 3093 3596
rect 3111 3576 3115 3596
rect 3121 3576 3125 3596
rect 3141 3556 3145 3596
rect 3205 3556 3209 3596
rect 3225 3556 3229 3596
rect 3245 3556 3249 3596
rect 3305 3576 3309 3596
rect 3351 3576 3355 3596
rect 3371 3576 3375 3596
rect 3431 3576 3435 3596
rect 3505 3576 3509 3596
rect 3525 3576 3529 3596
rect 3574 3556 3578 3596
rect 3582 3556 3586 3596
rect 3604 3576 3608 3596
rect 3671 3576 3675 3596
rect 3691 3576 3695 3596
rect 3711 3556 3715 3596
rect 3806 3556 3810 3596
rect 3814 3556 3818 3596
rect 3834 3556 3838 3596
rect 3842 3556 3846 3596
rect 3913 3556 3917 3596
rect 3923 3556 3927 3596
rect 3971 3556 3975 3596
rect 3993 3576 3997 3596
rect 4003 3576 4007 3596
rect 4023 3576 4027 3596
rect 4031 3576 4035 3596
rect 4077 3576 4081 3596
rect 4099 3576 4103 3596
rect 4109 3576 4113 3596
rect 4131 3576 4135 3596
rect 4141 3576 4145 3596
rect 4161 3556 4165 3596
rect 4211 3556 4215 3596
rect 4233 3576 4237 3596
rect 4243 3576 4247 3596
rect 4263 3576 4267 3596
rect 4271 3576 4275 3596
rect 4317 3576 4321 3596
rect 4339 3576 4343 3596
rect 4349 3576 4353 3596
rect 4371 3576 4375 3596
rect 4381 3576 4385 3596
rect 4401 3556 4405 3596
rect 4465 3556 4469 3596
rect 4485 3556 4489 3596
rect 4505 3556 4509 3596
rect 4525 3556 4529 3596
rect 4545 3556 4549 3596
rect 4565 3556 4569 3596
rect 4585 3556 4589 3596
rect 4605 3556 4609 3596
rect 4651 3556 4655 3596
rect 4671 3556 4675 3596
rect 4691 3556 4695 3596
rect 35 3144 39 3184
rect 55 3144 59 3164
rect 65 3144 69 3164
rect 87 3144 91 3164
rect 97 3144 101 3164
rect 119 3144 123 3164
rect 165 3144 169 3164
rect 173 3144 177 3164
rect 193 3144 197 3164
rect 203 3144 207 3164
rect 225 3144 229 3184
rect 306 3144 310 3184
rect 314 3144 318 3184
rect 334 3144 338 3184
rect 342 3144 346 3184
rect 413 3144 417 3184
rect 423 3144 427 3184
rect 471 3144 475 3184
rect 493 3144 497 3164
rect 503 3144 507 3164
rect 523 3144 527 3164
rect 531 3144 535 3164
rect 577 3144 581 3164
rect 599 3144 603 3164
rect 609 3144 613 3164
rect 631 3144 635 3164
rect 641 3144 645 3164
rect 661 3144 665 3184
rect 725 3144 729 3184
rect 745 3144 749 3184
rect 765 3144 769 3184
rect 846 3144 850 3184
rect 854 3144 858 3184
rect 874 3144 878 3184
rect 882 3144 886 3184
rect 933 3144 937 3184
rect 943 3144 947 3184
rect 1048 3144 1052 3204
rect 1056 3144 1060 3204
rect 1064 3144 1068 3204
rect 1135 3144 1139 3184
rect 1155 3144 1159 3184
rect 1165 3144 1169 3184
rect 1212 3144 1216 3204
rect 1220 3144 1224 3204
rect 1228 3144 1232 3204
rect 1311 3144 1315 3184
rect 1331 3144 1335 3184
rect 1351 3144 1355 3184
rect 1413 3144 1417 3184
rect 1423 3144 1427 3184
rect 1505 3144 1509 3184
rect 1525 3144 1529 3164
rect 1545 3144 1549 3164
rect 1613 3144 1617 3184
rect 1623 3144 1627 3184
rect 1671 3144 1675 3184
rect 1691 3144 1695 3184
rect 1711 3144 1715 3184
rect 1785 3144 1789 3184
rect 1805 3144 1809 3184
rect 1825 3144 1829 3184
rect 1873 3144 1877 3184
rect 1883 3144 1887 3184
rect 1951 3144 1955 3184
rect 1971 3144 1975 3184
rect 1991 3144 1995 3184
rect 2065 3144 2069 3184
rect 2085 3144 2089 3184
rect 2105 3144 2109 3184
rect 2151 3144 2155 3164
rect 2211 3144 2215 3184
rect 2231 3144 2235 3184
rect 2251 3144 2255 3184
rect 2325 3144 2329 3164
rect 2373 3144 2377 3184
rect 2383 3144 2387 3184
rect 2451 3144 2455 3184
rect 2473 3144 2477 3164
rect 2483 3144 2487 3164
rect 2503 3144 2507 3164
rect 2511 3144 2515 3164
rect 2557 3144 2561 3164
rect 2579 3144 2583 3164
rect 2589 3144 2593 3164
rect 2611 3144 2615 3164
rect 2621 3144 2625 3164
rect 2641 3144 2645 3184
rect 2691 3144 2695 3164
rect 2713 3144 2717 3184
rect 2771 3144 2775 3184
rect 2793 3144 2797 3164
rect 2803 3144 2807 3164
rect 2823 3144 2827 3164
rect 2831 3144 2835 3164
rect 2877 3144 2881 3164
rect 2899 3144 2903 3164
rect 2909 3144 2913 3164
rect 2931 3144 2935 3164
rect 2941 3144 2945 3164
rect 2961 3144 2965 3184
rect 3025 3144 3029 3184
rect 3045 3144 3049 3184
rect 3065 3144 3069 3184
rect 3125 3144 3129 3184
rect 3145 3144 3149 3184
rect 3165 3144 3169 3184
rect 3211 3144 3215 3184
rect 3231 3144 3235 3184
rect 3251 3144 3255 3184
rect 3325 3144 3329 3184
rect 3345 3144 3349 3184
rect 3365 3144 3369 3184
rect 3411 3144 3415 3184
rect 3431 3144 3435 3184
rect 3451 3144 3455 3184
rect 3513 3144 3517 3184
rect 3523 3144 3527 3184
rect 3593 3144 3597 3184
rect 3603 3144 3607 3184
rect 3673 3144 3677 3184
rect 3683 3144 3687 3184
rect 3753 3144 3757 3184
rect 3763 3144 3767 3184
rect 3831 3144 3835 3164
rect 3853 3144 3857 3184
rect 3933 3144 3937 3184
rect 3943 3144 3947 3184
rect 4005 3144 4009 3164
rect 4025 3144 4029 3164
rect 4071 3144 4075 3164
rect 4093 3144 4097 3184
rect 4165 3144 4169 3164
rect 4225 3144 4229 3184
rect 4245 3144 4249 3184
rect 4265 3144 4269 3184
rect 4325 3144 4329 3164
rect 4371 3144 4375 3184
rect 4391 3144 4395 3184
rect 4411 3144 4415 3184
rect 4493 3144 4497 3184
rect 4503 3144 4507 3184
rect 4555 3144 4559 3184
rect 4575 3144 4579 3164
rect 4585 3144 4589 3164
rect 4607 3144 4611 3164
rect 4617 3144 4621 3164
rect 4639 3144 4643 3164
rect 4685 3144 4689 3164
rect 4693 3144 4697 3164
rect 4713 3144 4717 3164
rect 4723 3144 4727 3164
rect 4745 3144 4749 3184
rect 66 3076 70 3116
rect 74 3076 78 3116
rect 94 3076 98 3116
rect 102 3076 106 3116
rect 175 3076 179 3116
rect 195 3076 199 3116
rect 205 3076 209 3116
rect 251 3076 255 3116
rect 273 3096 277 3116
rect 283 3096 287 3116
rect 303 3096 307 3116
rect 311 3096 315 3116
rect 357 3096 361 3116
rect 379 3096 383 3116
rect 389 3096 393 3116
rect 411 3096 415 3116
rect 421 3096 425 3116
rect 441 3076 445 3116
rect 491 3076 495 3116
rect 511 3076 515 3116
rect 531 3076 535 3116
rect 593 3076 597 3116
rect 603 3076 607 3116
rect 693 3076 697 3116
rect 703 3076 707 3116
rect 765 3096 769 3116
rect 785 3096 789 3116
rect 833 3076 837 3116
rect 843 3076 847 3116
rect 925 3076 929 3116
rect 945 3076 949 3116
rect 965 3076 969 3116
rect 1025 3076 1029 3116
rect 1045 3076 1049 3116
rect 1065 3076 1069 3116
rect 1125 3096 1129 3116
rect 1145 3096 1149 3116
rect 1205 3076 1209 3116
rect 1225 3076 1229 3116
rect 1245 3076 1249 3116
rect 1293 3076 1297 3116
rect 1303 3076 1307 3116
rect 1385 3076 1389 3116
rect 1433 3076 1437 3116
rect 1443 3076 1447 3116
rect 1513 3076 1517 3116
rect 1523 3076 1527 3116
rect 1591 3096 1595 3116
rect 1613 3076 1617 3116
rect 1671 3076 1675 3116
rect 1691 3076 1695 3116
rect 1711 3076 1715 3116
rect 1771 3076 1775 3116
rect 1791 3076 1795 3116
rect 1811 3076 1815 3116
rect 1871 3096 1875 3116
rect 1891 3096 1895 3116
rect 1954 3076 1958 3116
rect 1962 3076 1966 3116
rect 1984 3096 1988 3116
rect 2051 3096 2055 3116
rect 2111 3076 2115 3116
rect 2131 3076 2135 3116
rect 2151 3076 2155 3116
rect 2211 3096 2215 3116
rect 2231 3096 2235 3116
rect 2313 3076 2317 3116
rect 2323 3076 2327 3116
rect 2371 3076 2375 3116
rect 2391 3076 2395 3116
rect 2411 3076 2415 3116
rect 2471 3096 2475 3116
rect 2531 3076 2535 3116
rect 2551 3076 2555 3116
rect 2571 3076 2575 3116
rect 2631 3096 2635 3116
rect 2653 3076 2657 3116
rect 2713 3076 2717 3116
rect 2723 3076 2727 3116
rect 2795 3076 2799 3116
rect 2815 3096 2819 3116
rect 2825 3096 2829 3116
rect 2847 3096 2851 3116
rect 2857 3096 2861 3116
rect 2879 3096 2883 3116
rect 2925 3096 2929 3116
rect 2933 3096 2937 3116
rect 2953 3096 2957 3116
rect 2963 3096 2967 3116
rect 2985 3076 2989 3116
rect 3045 3096 3049 3116
rect 3065 3096 3069 3116
rect 3132 3096 3136 3116
rect 3154 3076 3158 3116
rect 3162 3076 3166 3116
rect 3211 3096 3215 3116
rect 3231 3096 3235 3116
rect 3295 3076 3299 3116
rect 3315 3096 3319 3116
rect 3325 3096 3329 3116
rect 3347 3096 3351 3116
rect 3357 3096 3361 3116
rect 3379 3096 3383 3116
rect 3425 3096 3429 3116
rect 3433 3096 3437 3116
rect 3453 3096 3457 3116
rect 3463 3096 3467 3116
rect 3485 3076 3489 3116
rect 3535 3076 3539 3116
rect 3555 3096 3559 3116
rect 3565 3096 3569 3116
rect 3587 3096 3591 3116
rect 3597 3096 3601 3116
rect 3619 3096 3623 3116
rect 3665 3096 3669 3116
rect 3673 3096 3677 3116
rect 3693 3096 3697 3116
rect 3703 3096 3707 3116
rect 3725 3076 3729 3116
rect 3771 3096 3775 3116
rect 3791 3096 3795 3116
rect 3865 3076 3869 3116
rect 3885 3076 3889 3116
rect 3905 3076 3909 3116
rect 3965 3076 3969 3116
rect 3985 3076 3989 3116
rect 4005 3076 4009 3116
rect 4051 3076 4055 3116
rect 4071 3076 4075 3116
rect 4091 3076 4095 3116
rect 4151 3076 4155 3116
rect 4171 3076 4175 3116
rect 4191 3076 4195 3116
rect 4251 3096 4255 3116
rect 4312 3056 4316 3116
rect 4320 3056 4324 3116
rect 4328 3056 4332 3116
rect 4411 3076 4415 3116
rect 4433 3096 4437 3116
rect 4443 3096 4447 3116
rect 4463 3096 4467 3116
rect 4471 3096 4475 3116
rect 4517 3096 4521 3116
rect 4539 3096 4543 3116
rect 4549 3096 4553 3116
rect 4571 3096 4575 3116
rect 4581 3096 4585 3116
rect 4601 3076 4605 3116
rect 4651 3076 4655 3116
rect 4671 3076 4675 3116
rect 4691 3076 4695 3116
rect 45 2664 49 2684
rect 105 2664 109 2704
rect 125 2664 129 2704
rect 145 2664 149 2704
rect 194 2664 198 2704
rect 202 2664 206 2704
rect 222 2664 226 2704
rect 230 2664 234 2704
rect 313 2664 317 2704
rect 323 2664 327 2704
rect 391 2664 395 2704
rect 401 2664 405 2704
rect 421 2664 425 2704
rect 505 2664 509 2704
rect 525 2664 529 2704
rect 545 2664 549 2704
rect 593 2664 597 2704
rect 603 2664 607 2704
rect 685 2664 689 2704
rect 745 2664 749 2704
rect 793 2664 797 2704
rect 803 2664 807 2704
rect 871 2664 875 2704
rect 881 2664 885 2704
rect 901 2664 905 2704
rect 985 2664 989 2704
rect 1005 2664 1009 2704
rect 1025 2664 1029 2704
rect 1073 2664 1077 2704
rect 1083 2664 1087 2704
rect 1165 2664 1169 2704
rect 1185 2664 1189 2704
rect 1205 2664 1209 2704
rect 1251 2664 1255 2704
rect 1273 2664 1277 2684
rect 1283 2664 1287 2684
rect 1303 2664 1307 2684
rect 1311 2664 1315 2684
rect 1357 2664 1361 2684
rect 1379 2664 1383 2684
rect 1389 2664 1393 2684
rect 1411 2664 1415 2684
rect 1421 2664 1425 2684
rect 1441 2664 1445 2704
rect 1503 2664 1507 2704
rect 1525 2664 1529 2684
rect 1575 2664 1579 2704
rect 1595 2664 1599 2684
rect 1605 2664 1609 2684
rect 1627 2664 1631 2684
rect 1637 2664 1641 2684
rect 1659 2664 1663 2684
rect 1705 2664 1709 2684
rect 1713 2664 1717 2684
rect 1733 2664 1737 2684
rect 1743 2664 1747 2684
rect 1765 2664 1769 2704
rect 1811 2664 1815 2704
rect 1831 2664 1835 2704
rect 1851 2664 1855 2704
rect 1911 2664 1915 2684
rect 1971 2664 1975 2704
rect 1991 2664 1995 2704
rect 2011 2664 2015 2704
rect 2031 2664 2035 2704
rect 2105 2664 2109 2684
rect 2125 2664 2129 2684
rect 2185 2664 2189 2684
rect 2205 2664 2209 2684
rect 2265 2664 2269 2684
rect 2285 2664 2289 2684
rect 2331 2664 2335 2684
rect 2405 2664 2409 2684
rect 2425 2664 2429 2684
rect 2471 2664 2475 2684
rect 2531 2664 2535 2704
rect 2541 2664 2545 2704
rect 2561 2664 2565 2704
rect 2631 2664 2635 2704
rect 2651 2664 2655 2704
rect 2671 2664 2675 2704
rect 2731 2664 2735 2704
rect 2751 2664 2755 2704
rect 2771 2664 2775 2704
rect 2833 2664 2837 2704
rect 2843 2664 2847 2704
rect 2915 2664 2919 2704
rect 2935 2664 2939 2684
rect 2945 2664 2949 2684
rect 2967 2664 2971 2684
rect 2977 2664 2981 2684
rect 2999 2664 3003 2684
rect 3045 2664 3049 2684
rect 3053 2664 3057 2684
rect 3073 2664 3077 2684
rect 3083 2664 3087 2684
rect 3105 2664 3109 2704
rect 3155 2664 3159 2704
rect 3175 2664 3179 2684
rect 3185 2664 3189 2684
rect 3207 2664 3211 2684
rect 3217 2664 3221 2684
rect 3239 2664 3243 2684
rect 3285 2664 3289 2684
rect 3293 2664 3297 2684
rect 3313 2664 3317 2684
rect 3323 2664 3327 2684
rect 3345 2664 3349 2704
rect 3405 2664 3409 2684
rect 3465 2664 3469 2684
rect 3485 2664 3489 2684
rect 3545 2664 3549 2704
rect 3595 2664 3599 2704
rect 3615 2664 3619 2684
rect 3625 2664 3629 2684
rect 3647 2664 3651 2684
rect 3657 2664 3661 2684
rect 3679 2664 3683 2684
rect 3725 2664 3729 2684
rect 3733 2664 3737 2684
rect 3753 2664 3757 2684
rect 3763 2664 3767 2684
rect 3785 2664 3789 2704
rect 3866 2664 3870 2704
rect 3874 2664 3878 2704
rect 3894 2664 3898 2704
rect 3902 2664 3906 2704
rect 3965 2664 3969 2684
rect 3985 2664 3989 2684
rect 4031 2664 4035 2704
rect 4051 2664 4055 2704
rect 4071 2664 4075 2704
rect 4145 2664 4149 2704
rect 4165 2664 4169 2704
rect 4185 2664 4189 2704
rect 4231 2664 4235 2684
rect 4251 2664 4255 2684
rect 4315 2664 4319 2704
rect 4335 2664 4339 2684
rect 4345 2664 4349 2684
rect 4367 2664 4371 2684
rect 4377 2664 4381 2684
rect 4399 2664 4403 2684
rect 4445 2664 4449 2684
rect 4453 2664 4457 2684
rect 4473 2664 4477 2684
rect 4483 2664 4487 2684
rect 4505 2664 4509 2704
rect 4551 2664 4555 2704
rect 4571 2664 4575 2704
rect 4591 2664 4595 2704
rect 4653 2664 4657 2704
rect 4663 2664 4667 2704
rect 32 2576 36 2636
rect 40 2576 44 2636
rect 48 2576 52 2636
rect 134 2596 138 2636
rect 142 2596 146 2636
rect 164 2616 168 2636
rect 245 2616 249 2636
rect 315 2596 319 2636
rect 335 2596 339 2636
rect 345 2596 349 2636
rect 412 2616 416 2636
rect 434 2596 438 2636
rect 442 2596 446 2636
rect 528 2576 532 2636
rect 536 2576 540 2636
rect 544 2576 548 2636
rect 605 2596 609 2636
rect 625 2596 629 2636
rect 645 2596 649 2636
rect 705 2596 709 2636
rect 773 2596 777 2636
rect 783 2596 787 2636
rect 868 2576 872 2636
rect 876 2576 880 2636
rect 884 2576 888 2636
rect 945 2596 949 2636
rect 965 2596 969 2636
rect 985 2596 989 2636
rect 1033 2596 1037 2636
rect 1043 2596 1047 2636
rect 1148 2576 1152 2636
rect 1156 2576 1160 2636
rect 1164 2576 1168 2636
rect 1225 2616 1229 2636
rect 1285 2596 1289 2636
rect 1305 2596 1309 2636
rect 1325 2596 1329 2636
rect 1373 2596 1377 2636
rect 1383 2596 1387 2636
rect 1451 2596 1455 2636
rect 1533 2596 1537 2636
rect 1543 2596 1547 2636
rect 1595 2596 1599 2636
rect 1615 2616 1619 2636
rect 1625 2616 1629 2636
rect 1647 2616 1651 2636
rect 1657 2616 1661 2636
rect 1679 2616 1683 2636
rect 1725 2616 1729 2636
rect 1733 2616 1737 2636
rect 1753 2616 1757 2636
rect 1763 2616 1767 2636
rect 1785 2596 1789 2636
rect 1833 2596 1837 2636
rect 1843 2596 1847 2636
rect 1913 2596 1917 2636
rect 1923 2596 1927 2636
rect 1992 2576 1996 2636
rect 2000 2576 2004 2636
rect 2008 2576 2012 2636
rect 2091 2616 2095 2636
rect 2111 2616 2115 2636
rect 2185 2616 2189 2636
rect 2245 2616 2249 2636
rect 2265 2616 2269 2636
rect 2325 2616 2329 2636
rect 2385 2596 2389 2636
rect 2405 2596 2409 2636
rect 2425 2596 2429 2636
rect 2471 2616 2475 2636
rect 2491 2616 2495 2636
rect 2551 2596 2555 2636
rect 2561 2596 2565 2636
rect 2581 2596 2585 2636
rect 2651 2596 2655 2636
rect 2671 2596 2675 2636
rect 2691 2596 2695 2636
rect 2773 2596 2777 2636
rect 2783 2596 2787 2636
rect 2831 2616 2835 2636
rect 2851 2616 2855 2636
rect 2871 2596 2875 2636
rect 2933 2596 2937 2636
rect 2943 2596 2947 2636
rect 3011 2616 3015 2636
rect 3033 2596 3037 2636
rect 3091 2596 3095 2636
rect 3111 2596 3115 2636
rect 3131 2596 3135 2636
rect 3203 2596 3207 2636
rect 3225 2616 3229 2636
rect 3293 2596 3297 2636
rect 3303 2596 3307 2636
rect 3354 2596 3358 2636
rect 3362 2596 3366 2636
rect 3382 2596 3386 2636
rect 3390 2596 3394 2636
rect 3471 2616 3475 2636
rect 3493 2596 3497 2636
rect 3563 2596 3567 2636
rect 3585 2616 3589 2636
rect 3635 2596 3639 2636
rect 3655 2616 3659 2636
rect 3665 2616 3669 2636
rect 3687 2616 3691 2636
rect 3697 2616 3701 2636
rect 3719 2616 3723 2636
rect 3765 2616 3769 2636
rect 3773 2616 3777 2636
rect 3793 2616 3797 2636
rect 3803 2616 3807 2636
rect 3825 2596 3829 2636
rect 3892 2616 3896 2636
rect 3914 2596 3918 2636
rect 3922 2596 3926 2636
rect 3971 2616 3975 2636
rect 3991 2616 3995 2636
rect 4051 2596 4055 2636
rect 4071 2596 4075 2636
rect 4091 2596 4095 2636
rect 4111 2596 4115 2636
rect 4131 2596 4135 2636
rect 4151 2596 4155 2636
rect 4171 2596 4175 2636
rect 4191 2596 4195 2636
rect 4255 2596 4259 2636
rect 4275 2616 4279 2636
rect 4285 2616 4289 2636
rect 4307 2616 4311 2636
rect 4317 2616 4321 2636
rect 4339 2616 4343 2636
rect 4385 2616 4389 2636
rect 4393 2616 4397 2636
rect 4413 2616 4417 2636
rect 4423 2616 4427 2636
rect 4445 2596 4449 2636
rect 4491 2596 4495 2636
rect 4511 2596 4515 2636
rect 4531 2596 4535 2636
rect 4593 2596 4597 2636
rect 4603 2596 4607 2636
rect 4673 2596 4677 2636
rect 4683 2596 4687 2636
rect 68 2184 72 2244
rect 76 2184 80 2244
rect 84 2184 88 2244
rect 145 2184 149 2224
rect 165 2184 169 2224
rect 185 2184 189 2224
rect 231 2184 235 2224
rect 251 2184 255 2224
rect 271 2184 275 2224
rect 332 2184 336 2244
rect 340 2184 344 2244
rect 348 2184 352 2244
rect 434 2184 438 2224
rect 442 2184 446 2224
rect 464 2184 468 2204
rect 531 2184 535 2224
rect 551 2184 555 2224
rect 571 2184 575 2224
rect 652 2184 656 2204
rect 674 2184 678 2224
rect 682 2184 686 2224
rect 731 2184 735 2204
rect 815 2184 819 2224
rect 835 2184 839 2224
rect 845 2184 849 2224
rect 893 2184 897 2224
rect 903 2184 907 2224
rect 971 2184 975 2224
rect 981 2184 985 2224
rect 1001 2184 1005 2224
rect 1085 2184 1089 2224
rect 1105 2184 1109 2224
rect 1125 2184 1129 2224
rect 1185 2184 1189 2224
rect 1205 2184 1209 2224
rect 1225 2184 1229 2224
rect 1275 2184 1279 2224
rect 1295 2184 1299 2204
rect 1305 2184 1309 2204
rect 1327 2184 1331 2204
rect 1337 2184 1341 2204
rect 1359 2184 1363 2204
rect 1405 2184 1409 2204
rect 1413 2184 1417 2204
rect 1433 2184 1437 2204
rect 1443 2184 1447 2204
rect 1465 2184 1469 2224
rect 1525 2184 1529 2224
rect 1545 2184 1549 2224
rect 1565 2184 1569 2224
rect 1615 2184 1619 2224
rect 1635 2184 1639 2204
rect 1645 2184 1649 2204
rect 1667 2184 1671 2204
rect 1677 2184 1681 2204
rect 1699 2184 1703 2204
rect 1745 2184 1749 2204
rect 1753 2184 1757 2204
rect 1773 2184 1777 2204
rect 1783 2184 1787 2204
rect 1805 2184 1809 2224
rect 1865 2184 1869 2204
rect 1925 2184 1929 2204
rect 1971 2184 1975 2224
rect 1991 2184 1995 2224
rect 2011 2184 2015 2224
rect 2075 2184 2079 2224
rect 2095 2184 2099 2204
rect 2105 2184 2109 2204
rect 2127 2184 2131 2204
rect 2137 2184 2141 2204
rect 2159 2184 2163 2204
rect 2205 2184 2209 2204
rect 2213 2184 2217 2204
rect 2233 2184 2237 2204
rect 2243 2184 2247 2204
rect 2265 2184 2269 2224
rect 2332 2184 2336 2204
rect 2354 2184 2358 2224
rect 2362 2184 2366 2224
rect 2432 2184 2436 2204
rect 2454 2184 2458 2224
rect 2462 2184 2466 2224
rect 2512 2184 2516 2244
rect 2520 2184 2524 2244
rect 2528 2184 2532 2244
rect 2611 2184 2615 2224
rect 2621 2184 2625 2224
rect 2641 2184 2645 2224
rect 2711 2184 2715 2224
rect 2733 2184 2737 2204
rect 2743 2184 2747 2204
rect 2763 2184 2767 2204
rect 2771 2184 2775 2204
rect 2817 2184 2821 2204
rect 2839 2184 2843 2204
rect 2849 2184 2853 2204
rect 2871 2184 2875 2204
rect 2881 2184 2885 2204
rect 2901 2184 2905 2224
rect 2965 2184 2969 2224
rect 2985 2184 2989 2224
rect 3005 2184 3009 2224
rect 3065 2184 3069 2224
rect 3085 2184 3089 2224
rect 3105 2184 3109 2224
rect 3151 2184 3155 2224
rect 3171 2184 3175 2224
rect 3191 2184 3195 2224
rect 3251 2184 3255 2224
rect 3273 2184 3277 2204
rect 3283 2184 3287 2204
rect 3303 2184 3307 2204
rect 3311 2184 3315 2204
rect 3357 2184 3361 2204
rect 3379 2184 3383 2204
rect 3389 2184 3393 2204
rect 3411 2184 3415 2204
rect 3421 2184 3425 2204
rect 3441 2184 3445 2224
rect 3505 2184 3509 2224
rect 3525 2184 3529 2224
rect 3545 2184 3549 2224
rect 3605 2184 3609 2204
rect 3625 2184 3629 2204
rect 3671 2184 3675 2204
rect 3691 2184 3695 2204
rect 3711 2184 3715 2224
rect 3793 2184 3797 2224
rect 3803 2184 3807 2224
rect 3886 2184 3890 2224
rect 3894 2184 3898 2224
rect 3914 2184 3918 2224
rect 3922 2184 3926 2224
rect 4006 2184 4010 2224
rect 4014 2184 4018 2224
rect 4034 2184 4038 2224
rect 4042 2184 4046 2224
rect 4095 2184 4099 2224
rect 4115 2184 4119 2204
rect 4125 2184 4129 2204
rect 4147 2184 4151 2204
rect 4157 2184 4161 2204
rect 4179 2184 4183 2204
rect 4225 2184 4229 2204
rect 4233 2184 4237 2204
rect 4253 2184 4257 2204
rect 4263 2184 4267 2204
rect 4285 2184 4289 2224
rect 4331 2184 4335 2224
rect 4353 2184 4357 2204
rect 4363 2184 4367 2204
rect 4383 2184 4387 2204
rect 4391 2184 4395 2204
rect 4437 2184 4441 2204
rect 4459 2184 4463 2204
rect 4469 2184 4473 2204
rect 4491 2184 4495 2204
rect 4501 2184 4505 2204
rect 4521 2184 4525 2224
rect 4571 2184 4575 2224
rect 4591 2184 4595 2224
rect 4611 2184 4615 2224
rect 4673 2184 4677 2224
rect 4683 2184 4687 2224
rect 43 2116 47 2156
rect 65 2136 69 2156
rect 125 2116 129 2156
rect 145 2116 149 2156
rect 165 2116 169 2156
rect 248 2096 252 2156
rect 256 2096 260 2156
rect 264 2096 268 2156
rect 314 2116 318 2156
rect 322 2116 326 2156
rect 344 2136 348 2156
rect 414 2116 418 2156
rect 422 2116 426 2156
rect 444 2136 448 2156
rect 512 2096 516 2156
rect 520 2096 524 2156
rect 528 2096 532 2156
rect 612 2096 616 2156
rect 620 2096 624 2156
rect 628 2096 632 2156
rect 714 2116 718 2156
rect 722 2116 726 2156
rect 744 2136 748 2156
rect 825 2116 829 2156
rect 845 2116 849 2156
rect 865 2116 869 2156
rect 912 2096 916 2156
rect 920 2096 924 2156
rect 928 2096 932 2156
rect 1012 2096 1016 2156
rect 1020 2096 1024 2156
rect 1028 2096 1032 2156
rect 1112 2096 1116 2156
rect 1120 2096 1124 2156
rect 1128 2096 1132 2156
rect 1214 2116 1218 2156
rect 1222 2116 1226 2156
rect 1244 2136 1248 2156
rect 1311 2136 1315 2156
rect 1331 2136 1335 2156
rect 1413 2116 1417 2156
rect 1423 2116 1427 2156
rect 1493 2116 1497 2156
rect 1503 2116 1507 2156
rect 1553 2116 1557 2156
rect 1563 2116 1567 2156
rect 1645 2116 1649 2156
rect 1665 2116 1669 2156
rect 1685 2116 1689 2156
rect 1734 2116 1738 2156
rect 1742 2116 1746 2156
rect 1764 2136 1768 2156
rect 1831 2136 1835 2156
rect 1851 2136 1855 2156
rect 1925 2116 1929 2156
rect 1945 2116 1949 2156
rect 1965 2116 1969 2156
rect 2011 2116 2015 2156
rect 2031 2116 2035 2156
rect 2051 2116 2055 2156
rect 2125 2116 2129 2156
rect 2145 2116 2149 2156
rect 2165 2116 2169 2156
rect 2225 2116 2229 2156
rect 2245 2116 2249 2156
rect 2265 2116 2269 2156
rect 2285 2116 2289 2156
rect 2305 2116 2309 2156
rect 2325 2116 2329 2156
rect 2345 2116 2349 2156
rect 2365 2116 2369 2156
rect 2413 2116 2417 2156
rect 2423 2116 2427 2156
rect 2515 2116 2519 2156
rect 2535 2116 2539 2156
rect 2545 2116 2549 2156
rect 2591 2136 2595 2156
rect 2611 2136 2615 2156
rect 2631 2116 2635 2156
rect 2713 2116 2717 2156
rect 2723 2116 2727 2156
rect 2773 2116 2777 2156
rect 2783 2116 2787 2156
rect 2855 2116 2859 2156
rect 2875 2136 2879 2156
rect 2885 2136 2889 2156
rect 2907 2136 2911 2156
rect 2917 2136 2921 2156
rect 2939 2136 2943 2156
rect 2985 2136 2989 2156
rect 2993 2136 2997 2156
rect 3013 2136 3017 2156
rect 3023 2136 3027 2156
rect 3045 2116 3049 2156
rect 3112 2136 3116 2156
rect 3134 2116 3138 2156
rect 3142 2116 3146 2156
rect 3191 2136 3195 2156
rect 3211 2136 3215 2156
rect 3306 2116 3310 2156
rect 3314 2116 3318 2156
rect 3334 2116 3338 2156
rect 3342 2116 3346 2156
rect 3395 2116 3399 2156
rect 3415 2136 3419 2156
rect 3425 2136 3429 2156
rect 3447 2136 3451 2156
rect 3457 2136 3461 2156
rect 3479 2136 3483 2156
rect 3525 2136 3529 2156
rect 3533 2136 3537 2156
rect 3553 2136 3557 2156
rect 3563 2136 3567 2156
rect 3585 2116 3589 2156
rect 3631 2116 3635 2156
rect 3651 2116 3655 2156
rect 3671 2116 3675 2156
rect 3735 2116 3739 2156
rect 3755 2136 3759 2156
rect 3765 2136 3769 2156
rect 3787 2136 3791 2156
rect 3797 2136 3801 2156
rect 3819 2136 3823 2156
rect 3865 2136 3869 2156
rect 3873 2136 3877 2156
rect 3893 2136 3897 2156
rect 3903 2136 3907 2156
rect 3925 2116 3929 2156
rect 3971 2116 3975 2156
rect 3993 2136 3997 2156
rect 4003 2136 4007 2156
rect 4023 2136 4027 2156
rect 4031 2136 4035 2156
rect 4077 2136 4081 2156
rect 4099 2136 4103 2156
rect 4109 2136 4113 2156
rect 4131 2136 4135 2156
rect 4141 2136 4145 2156
rect 4161 2116 4165 2156
rect 4246 2116 4250 2156
rect 4254 2116 4258 2156
rect 4274 2116 4278 2156
rect 4282 2116 4286 2156
rect 4331 2136 4335 2156
rect 4405 2136 4409 2156
rect 4425 2136 4429 2156
rect 4485 2136 4489 2156
rect 4505 2136 4509 2156
rect 4551 2116 4555 2156
rect 4573 2136 4577 2156
rect 4583 2136 4587 2156
rect 4603 2136 4607 2156
rect 4611 2136 4615 2156
rect 4657 2136 4661 2156
rect 4679 2136 4683 2156
rect 4689 2136 4693 2156
rect 4711 2136 4715 2156
rect 4721 2136 4725 2156
rect 4741 2116 4745 2156
rect 66 1704 70 1744
rect 74 1704 78 1744
rect 94 1704 98 1744
rect 102 1704 106 1744
rect 151 1704 155 1744
rect 171 1704 175 1744
rect 191 1704 195 1744
rect 253 1704 257 1744
rect 263 1704 267 1744
rect 368 1704 372 1764
rect 376 1704 380 1764
rect 384 1704 388 1764
rect 434 1704 438 1744
rect 442 1704 446 1744
rect 462 1704 466 1744
rect 470 1704 474 1744
rect 551 1704 555 1744
rect 561 1704 565 1744
rect 581 1704 585 1744
rect 665 1704 669 1744
rect 711 1704 715 1724
rect 733 1704 737 1744
rect 805 1704 809 1744
rect 825 1704 829 1744
rect 845 1704 849 1744
rect 891 1704 895 1744
rect 911 1704 915 1744
rect 931 1704 935 1744
rect 992 1704 996 1764
rect 1000 1704 1004 1764
rect 1008 1704 1012 1764
rect 1091 1704 1095 1724
rect 1152 1704 1156 1764
rect 1160 1704 1164 1764
rect 1168 1704 1172 1764
rect 1252 1704 1256 1764
rect 1260 1704 1264 1764
rect 1268 1704 1272 1764
rect 1365 1704 1369 1724
rect 1446 1704 1450 1744
rect 1454 1704 1458 1744
rect 1474 1704 1478 1744
rect 1482 1704 1486 1744
rect 1532 1704 1536 1764
rect 1540 1704 1544 1764
rect 1548 1704 1552 1764
rect 1631 1704 1635 1724
rect 1705 1704 1709 1744
rect 1788 1704 1792 1764
rect 1796 1704 1800 1764
rect 1804 1704 1808 1764
rect 1851 1704 1855 1744
rect 1861 1704 1865 1744
rect 1881 1704 1885 1744
rect 1955 1704 1959 1744
rect 1975 1704 1979 1724
rect 1985 1704 1989 1724
rect 2007 1704 2011 1724
rect 2017 1704 2021 1724
rect 2039 1704 2043 1724
rect 2085 1704 2089 1724
rect 2093 1704 2097 1724
rect 2113 1704 2117 1724
rect 2123 1704 2127 1724
rect 2145 1704 2149 1744
rect 2205 1704 2209 1724
rect 2225 1704 2229 1724
rect 2271 1704 2275 1724
rect 2331 1704 2335 1744
rect 2351 1704 2355 1744
rect 2371 1704 2375 1744
rect 2431 1704 2435 1724
rect 2451 1704 2455 1724
rect 2511 1704 2515 1724
rect 2531 1704 2535 1724
rect 2591 1704 2595 1744
rect 2611 1704 2615 1744
rect 2631 1704 2635 1744
rect 2713 1704 2717 1744
rect 2723 1704 2727 1744
rect 2785 1704 2789 1724
rect 2805 1704 2809 1724
rect 2851 1704 2855 1744
rect 2871 1704 2875 1744
rect 2891 1704 2895 1744
rect 2951 1704 2955 1724
rect 3025 1704 3029 1724
rect 3045 1704 3049 1724
rect 3091 1704 3095 1744
rect 3113 1704 3117 1724
rect 3123 1704 3127 1724
rect 3143 1704 3147 1724
rect 3151 1704 3155 1724
rect 3197 1704 3201 1724
rect 3219 1704 3223 1724
rect 3229 1704 3233 1724
rect 3251 1704 3255 1724
rect 3261 1704 3265 1724
rect 3281 1704 3285 1744
rect 3331 1704 3335 1744
rect 3351 1704 3355 1744
rect 3371 1704 3375 1744
rect 3433 1704 3437 1744
rect 3443 1704 3447 1744
rect 3511 1704 3515 1744
rect 3533 1704 3537 1724
rect 3543 1704 3547 1724
rect 3563 1704 3567 1724
rect 3571 1704 3575 1724
rect 3617 1704 3621 1724
rect 3639 1704 3643 1724
rect 3649 1704 3653 1724
rect 3671 1704 3675 1724
rect 3681 1704 3685 1724
rect 3701 1704 3705 1744
rect 3751 1704 3755 1724
rect 3773 1704 3777 1744
rect 3853 1704 3857 1744
rect 3863 1704 3867 1744
rect 3925 1704 3929 1744
rect 3945 1704 3949 1744
rect 3965 1704 3969 1744
rect 4025 1704 4029 1744
rect 4045 1704 4049 1744
rect 4065 1704 4069 1744
rect 4111 1704 4115 1724
rect 4131 1704 4135 1724
rect 4151 1704 4155 1744
rect 4225 1704 4229 1724
rect 4274 1704 4278 1744
rect 4282 1704 4286 1744
rect 4304 1704 4308 1724
rect 4385 1704 4389 1724
rect 4405 1704 4409 1724
rect 4451 1704 4455 1744
rect 4473 1704 4477 1724
rect 4483 1704 4487 1724
rect 4503 1704 4507 1724
rect 4511 1704 4515 1724
rect 4557 1704 4561 1724
rect 4579 1704 4583 1724
rect 4589 1704 4593 1724
rect 4611 1704 4615 1724
rect 4621 1704 4625 1724
rect 4641 1704 4645 1744
rect 4713 1704 4717 1744
rect 4723 1704 4727 1744
rect 45 1656 49 1676
rect 112 1656 116 1676
rect 134 1636 138 1676
rect 142 1636 146 1676
rect 192 1616 196 1676
rect 200 1616 204 1676
rect 208 1616 212 1676
rect 293 1636 297 1676
rect 303 1636 307 1676
rect 385 1636 389 1676
rect 405 1636 409 1676
rect 425 1636 429 1676
rect 483 1636 487 1676
rect 505 1656 509 1676
rect 565 1656 569 1676
rect 612 1616 616 1676
rect 620 1616 624 1676
rect 628 1616 632 1676
rect 714 1636 718 1676
rect 722 1636 726 1676
rect 744 1656 748 1676
rect 812 1616 816 1676
rect 820 1616 824 1676
rect 828 1616 832 1676
rect 914 1636 918 1676
rect 922 1636 926 1676
rect 944 1656 948 1676
rect 1012 1616 1016 1676
rect 1020 1616 1024 1676
rect 1028 1616 1032 1676
rect 1125 1636 1129 1676
rect 1145 1636 1149 1676
rect 1165 1636 1169 1676
rect 1212 1616 1216 1676
rect 1220 1616 1224 1676
rect 1228 1616 1232 1676
rect 1314 1636 1318 1676
rect 1322 1636 1326 1676
rect 1344 1656 1348 1676
rect 1425 1656 1429 1676
rect 1472 1616 1476 1676
rect 1480 1616 1484 1676
rect 1488 1616 1492 1676
rect 1574 1636 1578 1676
rect 1582 1636 1586 1676
rect 1604 1656 1608 1676
rect 1672 1616 1676 1676
rect 1680 1616 1684 1676
rect 1688 1616 1692 1676
rect 1771 1636 1775 1676
rect 1791 1636 1795 1676
rect 1811 1636 1815 1676
rect 1892 1656 1896 1676
rect 1914 1636 1918 1676
rect 1922 1636 1926 1676
rect 1971 1656 1975 1676
rect 2032 1616 2036 1676
rect 2040 1616 2044 1676
rect 2048 1616 2052 1676
rect 2145 1636 2149 1676
rect 2165 1636 2169 1676
rect 2185 1636 2189 1676
rect 2231 1656 2235 1676
rect 2291 1636 2295 1676
rect 2313 1656 2317 1676
rect 2323 1656 2327 1676
rect 2343 1656 2347 1676
rect 2351 1656 2355 1676
rect 2397 1656 2401 1676
rect 2419 1656 2423 1676
rect 2429 1656 2433 1676
rect 2451 1656 2455 1676
rect 2461 1656 2465 1676
rect 2481 1636 2485 1676
rect 2545 1636 2549 1676
rect 2565 1636 2569 1676
rect 2585 1636 2589 1676
rect 2655 1636 2659 1676
rect 2675 1636 2679 1676
rect 2685 1636 2689 1676
rect 2731 1656 2735 1676
rect 2751 1656 2755 1676
rect 2814 1636 2818 1676
rect 2822 1636 2826 1676
rect 2844 1656 2848 1676
rect 2925 1656 2929 1676
rect 2945 1656 2949 1676
rect 3005 1656 3009 1676
rect 3065 1656 3069 1676
rect 3111 1636 3115 1676
rect 3131 1636 3135 1676
rect 3151 1636 3155 1676
rect 3213 1636 3217 1676
rect 3223 1636 3227 1676
rect 3313 1636 3317 1676
rect 3323 1636 3327 1676
rect 3385 1636 3389 1676
rect 3405 1636 3409 1676
rect 3425 1636 3429 1676
rect 3475 1636 3479 1676
rect 3495 1656 3499 1676
rect 3505 1656 3509 1676
rect 3527 1656 3531 1676
rect 3537 1656 3541 1676
rect 3559 1656 3563 1676
rect 3605 1656 3609 1676
rect 3613 1656 3617 1676
rect 3633 1656 3637 1676
rect 3643 1656 3647 1676
rect 3665 1636 3669 1676
rect 3711 1656 3715 1676
rect 3785 1656 3789 1676
rect 3845 1636 3849 1676
rect 3865 1636 3869 1676
rect 3885 1636 3889 1676
rect 3931 1656 3935 1676
rect 3951 1656 3955 1676
rect 4011 1656 4015 1676
rect 4031 1656 4035 1676
rect 4091 1656 4095 1676
rect 4154 1636 4158 1676
rect 4162 1636 4166 1676
rect 4184 1656 4188 1676
rect 4251 1656 4255 1676
rect 4271 1656 4275 1676
rect 4334 1636 4338 1676
rect 4342 1636 4346 1676
rect 4364 1656 4368 1676
rect 4431 1656 4435 1676
rect 4491 1656 4495 1676
rect 4565 1656 4569 1676
rect 4611 1636 4615 1676
rect 4631 1636 4635 1676
rect 4651 1636 4655 1676
rect 4713 1636 4717 1676
rect 4723 1636 4727 1676
rect 52 1224 56 1244
rect 74 1224 78 1264
rect 82 1224 86 1264
rect 132 1224 136 1284
rect 140 1224 144 1284
rect 148 1224 152 1284
rect 232 1224 236 1284
rect 240 1224 244 1284
rect 248 1224 252 1284
rect 353 1224 357 1264
rect 363 1224 367 1264
rect 411 1224 415 1264
rect 431 1224 435 1264
rect 451 1224 455 1264
rect 514 1224 518 1264
rect 522 1224 526 1264
rect 544 1224 548 1244
rect 611 1224 615 1264
rect 631 1224 635 1264
rect 651 1224 655 1264
rect 711 1224 715 1264
rect 731 1224 735 1264
rect 751 1224 755 1264
rect 811 1224 815 1264
rect 821 1224 825 1264
rect 841 1224 845 1264
rect 933 1224 937 1264
rect 943 1224 947 1264
rect 993 1224 997 1264
rect 1003 1224 1007 1264
rect 1108 1224 1112 1284
rect 1116 1224 1120 1284
rect 1124 1224 1128 1284
rect 1185 1224 1189 1244
rect 1255 1224 1259 1264
rect 1275 1224 1279 1264
rect 1285 1224 1289 1264
rect 1331 1224 1335 1264
rect 1351 1224 1355 1264
rect 1371 1224 1375 1264
rect 1445 1224 1449 1264
rect 1465 1224 1469 1264
rect 1485 1224 1489 1264
rect 1533 1224 1537 1264
rect 1543 1224 1547 1264
rect 1611 1224 1615 1264
rect 1631 1224 1635 1264
rect 1651 1224 1655 1264
rect 1713 1224 1717 1264
rect 1723 1224 1727 1264
rect 1794 1224 1798 1264
rect 1802 1224 1806 1264
rect 1824 1224 1828 1244
rect 1892 1224 1896 1284
rect 1900 1224 1904 1284
rect 1908 1224 1912 1284
rect 1991 1224 1995 1264
rect 2011 1224 2015 1264
rect 2031 1224 2035 1264
rect 2091 1224 2095 1244
rect 2152 1224 2156 1284
rect 2160 1224 2164 1284
rect 2168 1224 2172 1284
rect 2253 1224 2257 1264
rect 2263 1224 2267 1264
rect 2331 1224 2335 1244
rect 2351 1224 2355 1244
rect 2371 1224 2375 1264
rect 2453 1224 2457 1264
rect 2463 1224 2467 1264
rect 2511 1224 2515 1244
rect 2583 1224 2587 1264
rect 2605 1224 2609 1244
rect 2651 1224 2655 1264
rect 2671 1224 2675 1264
rect 2691 1224 2695 1264
rect 2765 1224 2769 1264
rect 2785 1224 2789 1264
rect 2805 1224 2809 1264
rect 2825 1224 2829 1264
rect 2875 1224 2879 1264
rect 2895 1224 2899 1244
rect 2905 1224 2909 1244
rect 2927 1224 2931 1244
rect 2937 1224 2941 1244
rect 2959 1224 2963 1244
rect 3005 1224 3009 1244
rect 3013 1224 3017 1244
rect 3033 1224 3037 1244
rect 3043 1224 3047 1244
rect 3065 1224 3069 1264
rect 3125 1224 3129 1244
rect 3145 1224 3149 1244
rect 3212 1224 3216 1244
rect 3234 1224 3238 1264
rect 3242 1224 3246 1264
rect 3295 1224 3299 1264
rect 3315 1224 3319 1244
rect 3325 1224 3329 1244
rect 3347 1224 3351 1244
rect 3357 1224 3361 1244
rect 3379 1224 3383 1244
rect 3425 1224 3429 1244
rect 3433 1224 3437 1244
rect 3453 1224 3457 1244
rect 3463 1224 3467 1244
rect 3485 1224 3489 1264
rect 3545 1224 3549 1244
rect 3605 1224 3609 1244
rect 3625 1224 3629 1244
rect 3685 1224 3689 1244
rect 3705 1224 3709 1244
rect 3751 1224 3755 1244
rect 3811 1224 3815 1264
rect 3833 1224 3837 1244
rect 3843 1224 3847 1244
rect 3863 1224 3867 1244
rect 3871 1224 3875 1244
rect 3917 1224 3921 1244
rect 3939 1224 3943 1244
rect 3949 1224 3953 1244
rect 3971 1224 3975 1244
rect 3981 1224 3985 1244
rect 4001 1224 4005 1264
rect 4051 1224 4055 1264
rect 4071 1224 4075 1264
rect 4091 1224 4095 1264
rect 4153 1224 4157 1264
rect 4163 1224 4167 1264
rect 4243 1224 4247 1264
rect 4265 1224 4269 1244
rect 4333 1224 4337 1264
rect 4343 1224 4347 1264
rect 4405 1224 4409 1264
rect 4425 1224 4429 1264
rect 4445 1224 4449 1264
rect 4505 1224 4509 1264
rect 4525 1224 4529 1264
rect 4545 1224 4549 1264
rect 4591 1224 4595 1244
rect 4611 1224 4615 1244
rect 4671 1224 4675 1244
rect 4745 1224 4749 1244
rect 45 1156 49 1196
rect 65 1156 69 1196
rect 85 1156 89 1196
rect 131 1156 135 1196
rect 151 1156 155 1196
rect 171 1156 175 1196
rect 232 1136 236 1196
rect 240 1136 244 1196
rect 248 1136 252 1196
rect 334 1156 338 1196
rect 342 1156 346 1196
rect 364 1176 368 1196
rect 432 1136 436 1196
rect 440 1136 444 1196
rect 448 1136 452 1196
rect 534 1156 538 1196
rect 542 1156 546 1196
rect 564 1176 568 1196
rect 653 1156 657 1196
rect 663 1156 667 1196
rect 735 1156 739 1196
rect 755 1156 759 1196
rect 765 1156 769 1196
rect 848 1136 852 1196
rect 856 1136 860 1196
rect 864 1136 868 1196
rect 925 1156 929 1196
rect 945 1156 949 1196
rect 965 1156 969 1196
rect 1011 1156 1015 1196
rect 1031 1156 1035 1196
rect 1051 1156 1055 1196
rect 1125 1156 1129 1196
rect 1145 1156 1149 1196
rect 1165 1156 1169 1196
rect 1233 1156 1237 1196
rect 1243 1156 1247 1196
rect 1315 1156 1319 1196
rect 1335 1156 1339 1196
rect 1345 1156 1349 1196
rect 1393 1156 1397 1196
rect 1403 1156 1407 1196
rect 1485 1156 1489 1196
rect 1553 1156 1557 1196
rect 1563 1156 1567 1196
rect 1633 1156 1637 1196
rect 1643 1156 1647 1196
rect 1692 1136 1696 1196
rect 1700 1136 1704 1196
rect 1708 1136 1712 1196
rect 1813 1156 1817 1196
rect 1823 1156 1827 1196
rect 1872 1136 1876 1196
rect 1880 1136 1884 1196
rect 1888 1136 1892 1196
rect 1973 1156 1977 1196
rect 1983 1156 1987 1196
rect 2086 1156 2090 1196
rect 2094 1156 2098 1196
rect 2114 1156 2118 1196
rect 2122 1156 2126 1196
rect 2208 1136 2212 1196
rect 2216 1136 2220 1196
rect 2224 1136 2228 1196
rect 2293 1156 2297 1196
rect 2303 1156 2307 1196
rect 2354 1156 2358 1196
rect 2362 1156 2366 1196
rect 2384 1176 2388 1196
rect 2465 1176 2469 1196
rect 2533 1156 2537 1196
rect 2543 1156 2547 1196
rect 2605 1156 2609 1196
rect 2625 1156 2629 1196
rect 2645 1156 2649 1196
rect 2665 1156 2669 1196
rect 2711 1176 2715 1196
rect 2733 1156 2737 1196
rect 2795 1156 2799 1196
rect 2815 1176 2819 1196
rect 2825 1176 2829 1196
rect 2847 1176 2851 1196
rect 2857 1176 2861 1196
rect 2879 1176 2883 1196
rect 2925 1176 2929 1196
rect 2933 1176 2937 1196
rect 2953 1176 2957 1196
rect 2963 1176 2967 1196
rect 2985 1156 2989 1196
rect 3033 1156 3037 1196
rect 3043 1156 3047 1196
rect 3125 1156 3129 1196
rect 3145 1156 3149 1196
rect 3165 1156 3169 1196
rect 3211 1156 3215 1196
rect 3231 1156 3235 1196
rect 3251 1156 3255 1196
rect 3271 1156 3275 1196
rect 3343 1156 3347 1196
rect 3365 1176 3369 1196
rect 3411 1176 3415 1196
rect 3433 1156 3437 1196
rect 3491 1156 3495 1196
rect 3511 1156 3515 1196
rect 3531 1156 3535 1196
rect 3551 1156 3555 1196
rect 3571 1156 3575 1196
rect 3591 1156 3595 1196
rect 3611 1156 3615 1196
rect 3631 1156 3635 1196
rect 3691 1156 3695 1196
rect 3711 1156 3715 1196
rect 3731 1156 3735 1196
rect 3751 1156 3755 1196
rect 3771 1156 3775 1196
rect 3791 1156 3795 1196
rect 3811 1156 3815 1196
rect 3831 1156 3835 1196
rect 3891 1176 3895 1196
rect 3913 1156 3917 1196
rect 3973 1156 3977 1196
rect 3983 1156 3987 1196
rect 4051 1156 4055 1196
rect 4073 1176 4077 1196
rect 4083 1176 4087 1196
rect 4103 1176 4107 1196
rect 4111 1176 4115 1196
rect 4157 1176 4161 1196
rect 4179 1176 4183 1196
rect 4189 1176 4193 1196
rect 4211 1176 4215 1196
rect 4221 1176 4225 1196
rect 4241 1156 4245 1196
rect 4293 1156 4297 1196
rect 4303 1156 4307 1196
rect 4371 1156 4375 1196
rect 4391 1156 4395 1196
rect 4411 1156 4415 1196
rect 4493 1156 4497 1196
rect 4503 1156 4507 1196
rect 4551 1156 4555 1196
rect 4571 1156 4575 1196
rect 4591 1156 4595 1196
rect 4652 1136 4656 1196
rect 4660 1136 4664 1196
rect 4668 1136 4672 1196
rect 53 744 57 784
rect 63 744 67 784
rect 135 744 139 784
rect 155 744 159 784
rect 165 744 169 784
rect 225 744 229 784
rect 245 744 249 784
rect 265 744 269 784
rect 346 744 350 784
rect 354 744 358 784
rect 374 744 378 784
rect 382 744 386 784
rect 443 744 447 784
rect 465 744 469 764
rect 511 744 515 764
rect 585 744 589 764
rect 652 744 656 764
rect 674 744 678 784
rect 682 744 686 784
rect 732 744 736 804
rect 740 744 744 804
rect 748 744 752 804
rect 855 744 859 784
rect 875 744 879 784
rect 885 744 889 784
rect 933 744 937 784
rect 943 744 947 784
rect 1048 744 1052 804
rect 1056 744 1060 804
rect 1064 744 1068 804
rect 1111 744 1115 784
rect 1131 744 1135 784
rect 1151 744 1155 784
rect 1248 744 1252 804
rect 1256 744 1260 804
rect 1264 744 1268 804
rect 1311 744 1315 764
rect 1371 744 1375 784
rect 1391 744 1395 784
rect 1411 744 1415 784
rect 1493 744 1497 784
rect 1503 744 1507 784
rect 1553 744 1557 784
rect 1563 744 1567 784
rect 1645 744 1649 784
rect 1665 744 1669 784
rect 1685 744 1689 784
rect 1731 744 1735 784
rect 1741 744 1745 784
rect 1761 744 1765 784
rect 1845 744 1849 764
rect 1913 744 1917 784
rect 1923 744 1927 784
rect 1971 744 1975 764
rect 2068 744 2072 804
rect 2076 744 2080 804
rect 2084 744 2088 804
rect 2131 744 2135 764
rect 2191 744 2195 784
rect 2211 744 2215 784
rect 2231 744 2235 784
rect 2312 744 2316 764
rect 2334 744 2338 784
rect 2342 744 2346 784
rect 2391 744 2395 764
rect 2452 744 2456 804
rect 2460 744 2464 804
rect 2468 744 2472 804
rect 2588 744 2592 804
rect 2596 744 2600 804
rect 2604 744 2608 804
rect 2654 744 2658 784
rect 2662 744 2666 784
rect 2684 744 2688 764
rect 2773 744 2777 784
rect 2783 744 2787 784
rect 2845 744 2849 784
rect 2865 744 2869 784
rect 2885 744 2889 784
rect 2905 744 2909 784
rect 2965 744 2969 764
rect 3025 744 3029 764
rect 3045 744 3049 764
rect 3105 744 3109 764
rect 3125 744 3129 764
rect 3171 744 3175 764
rect 3231 744 3235 784
rect 3251 744 3255 784
rect 3271 744 3275 784
rect 3333 744 3337 784
rect 3343 744 3347 784
rect 3411 744 3415 784
rect 3433 744 3437 764
rect 3443 744 3447 764
rect 3463 744 3467 764
rect 3471 744 3475 764
rect 3517 744 3521 764
rect 3539 744 3543 764
rect 3549 744 3553 764
rect 3571 744 3575 764
rect 3581 744 3585 764
rect 3601 744 3605 784
rect 3651 744 3655 764
rect 3673 744 3677 784
rect 3735 744 3739 784
rect 3755 744 3759 764
rect 3765 744 3769 764
rect 3787 744 3791 764
rect 3797 744 3801 764
rect 3819 744 3823 764
rect 3865 744 3869 764
rect 3873 744 3877 764
rect 3893 744 3897 764
rect 3903 744 3907 764
rect 3925 744 3929 784
rect 3985 744 3989 784
rect 4005 744 4009 784
rect 4025 744 4029 784
rect 4071 744 4075 784
rect 4093 744 4097 764
rect 4103 744 4107 764
rect 4123 744 4127 764
rect 4131 744 4135 764
rect 4177 744 4181 764
rect 4199 744 4203 764
rect 4209 744 4213 764
rect 4231 744 4235 764
rect 4241 744 4245 764
rect 4261 744 4265 784
rect 4315 744 4319 784
rect 4335 744 4339 764
rect 4345 744 4349 764
rect 4367 744 4371 764
rect 4377 744 4381 764
rect 4399 744 4403 764
rect 4445 744 4449 764
rect 4453 744 4457 764
rect 4473 744 4477 764
rect 4483 744 4487 764
rect 4505 744 4509 784
rect 4551 744 4555 784
rect 4571 744 4575 784
rect 4591 744 4595 784
rect 4651 744 4655 784
rect 4671 744 4675 784
rect 4691 744 4695 784
rect 45 696 49 716
rect 65 696 69 716
rect 132 696 136 716
rect 154 676 158 716
rect 162 676 166 716
rect 211 696 215 716
rect 292 696 296 716
rect 314 676 318 716
rect 322 676 326 716
rect 372 656 376 716
rect 380 656 384 716
rect 388 656 392 716
rect 485 676 489 716
rect 505 676 509 716
rect 525 676 529 716
rect 583 676 587 716
rect 605 696 609 716
rect 665 676 669 716
rect 685 676 689 716
rect 705 676 709 716
rect 763 676 767 716
rect 785 696 789 716
rect 831 676 835 716
rect 841 676 845 716
rect 861 676 865 716
rect 931 676 935 716
rect 951 676 955 716
rect 971 676 975 716
rect 1045 676 1049 716
rect 1065 676 1069 716
rect 1085 676 1089 716
rect 1145 676 1149 716
rect 1194 676 1198 716
rect 1202 676 1206 716
rect 1224 696 1228 716
rect 1305 696 1309 716
rect 1351 676 1355 716
rect 1371 676 1375 716
rect 1391 676 1395 716
rect 1451 676 1455 716
rect 1471 676 1475 716
rect 1491 676 1495 716
rect 1572 696 1576 716
rect 1594 676 1598 716
rect 1602 676 1606 716
rect 1654 676 1658 716
rect 1662 676 1666 716
rect 1684 696 1688 716
rect 1752 656 1756 716
rect 1760 656 1764 716
rect 1768 656 1772 716
rect 1851 676 1855 716
rect 1871 676 1875 716
rect 1891 676 1895 716
rect 1972 696 1976 716
rect 1994 676 1998 716
rect 2002 676 2006 716
rect 2051 676 2055 716
rect 2071 676 2075 716
rect 2091 676 2095 716
rect 2188 656 2192 716
rect 2196 656 2200 716
rect 2204 656 2208 716
rect 2265 676 2269 716
rect 2285 676 2289 716
rect 2305 676 2309 716
rect 2351 676 2355 716
rect 2371 676 2375 716
rect 2391 676 2395 716
rect 2452 656 2456 716
rect 2460 656 2464 716
rect 2468 656 2472 716
rect 2552 656 2556 716
rect 2560 656 2564 716
rect 2568 656 2572 716
rect 2665 696 2669 716
rect 2712 656 2716 716
rect 2720 656 2724 716
rect 2728 656 2732 716
rect 2815 676 2819 716
rect 2835 696 2839 716
rect 2845 696 2849 716
rect 2867 696 2871 716
rect 2877 696 2881 716
rect 2899 696 2903 716
rect 2945 696 2949 716
rect 2953 696 2957 716
rect 2973 696 2977 716
rect 2983 696 2987 716
rect 3005 676 3009 716
rect 3051 676 3055 716
rect 3071 676 3075 716
rect 3091 676 3095 716
rect 3151 696 3155 716
rect 3211 696 3215 716
rect 3272 656 3276 716
rect 3280 656 3284 716
rect 3288 656 3292 716
rect 3385 696 3389 716
rect 3453 676 3457 716
rect 3463 676 3467 716
rect 3525 676 3529 716
rect 3545 676 3549 716
rect 3565 676 3569 716
rect 3615 676 3619 716
rect 3635 696 3639 716
rect 3645 696 3649 716
rect 3667 696 3671 716
rect 3677 696 3681 716
rect 3699 696 3703 716
rect 3745 696 3749 716
rect 3753 696 3757 716
rect 3773 696 3777 716
rect 3783 696 3787 716
rect 3805 676 3809 716
rect 3851 676 3855 716
rect 3871 676 3875 716
rect 3891 676 3895 716
rect 3973 676 3977 716
rect 3983 676 3987 716
rect 4031 676 4035 716
rect 4053 696 4057 716
rect 4063 696 4067 716
rect 4083 696 4087 716
rect 4091 696 4095 716
rect 4137 696 4141 716
rect 4159 696 4163 716
rect 4169 696 4173 716
rect 4191 696 4195 716
rect 4201 696 4205 716
rect 4221 676 4225 716
rect 4273 676 4277 716
rect 4283 676 4287 716
rect 4353 676 4357 716
rect 4363 676 4367 716
rect 4445 676 4449 716
rect 4465 676 4469 716
rect 4485 676 4489 716
rect 4535 676 4539 716
rect 4555 696 4559 716
rect 4565 696 4569 716
rect 4587 696 4591 716
rect 4597 696 4601 716
rect 4619 696 4623 716
rect 4665 696 4669 716
rect 4673 696 4677 716
rect 4693 696 4697 716
rect 4703 696 4707 716
rect 4725 676 4729 716
rect 33 264 37 304
rect 43 264 47 304
rect 113 264 117 304
rect 123 264 127 304
rect 213 264 217 304
rect 223 264 227 304
rect 293 264 297 304
rect 303 264 307 304
rect 375 264 379 304
rect 395 264 399 304
rect 405 264 409 304
rect 473 264 477 304
rect 483 264 487 304
rect 568 264 572 324
rect 576 264 580 324
rect 584 264 588 324
rect 666 264 670 304
rect 674 264 678 304
rect 694 264 698 304
rect 702 264 706 304
rect 765 264 769 284
rect 785 264 789 284
rect 853 264 857 304
rect 863 264 867 304
rect 913 264 917 304
rect 923 264 927 304
rect 1013 264 1017 304
rect 1023 264 1027 304
rect 1093 264 1097 304
rect 1103 264 1107 304
rect 1186 264 1190 304
rect 1194 264 1198 304
rect 1214 264 1218 304
rect 1222 264 1226 304
rect 1271 264 1275 304
rect 1291 264 1295 304
rect 1311 264 1315 304
rect 1385 264 1389 284
rect 1405 264 1409 284
rect 1451 264 1455 304
rect 1471 264 1475 304
rect 1491 264 1495 304
rect 1551 264 1555 284
rect 1632 264 1636 284
rect 1654 264 1658 304
rect 1662 264 1666 304
rect 1711 264 1715 284
rect 1772 264 1776 324
rect 1780 264 1784 324
rect 1788 264 1792 324
rect 1874 264 1878 304
rect 1882 264 1886 304
rect 1904 264 1908 284
rect 1973 264 1977 304
rect 1983 264 1987 304
rect 2053 264 2057 304
rect 2063 264 2067 304
rect 2133 264 2137 304
rect 2143 264 2147 304
rect 2225 264 2229 284
rect 2245 264 2249 284
rect 2313 264 2317 304
rect 2323 264 2327 304
rect 2371 264 2375 284
rect 2391 264 2395 284
rect 2452 264 2456 324
rect 2460 264 2464 324
rect 2468 264 2472 324
rect 2565 264 2569 284
rect 2648 264 2652 324
rect 2656 264 2660 324
rect 2664 264 2668 324
rect 2714 264 2718 304
rect 2722 264 2726 304
rect 2744 264 2748 284
rect 2811 264 2815 284
rect 2831 264 2835 284
rect 2913 264 2917 304
rect 2923 264 2927 304
rect 2985 264 2989 304
rect 3005 264 3009 304
rect 3025 264 3029 304
rect 3085 264 3089 304
rect 3105 264 3109 304
rect 3125 264 3129 304
rect 3185 264 3189 284
rect 3205 264 3209 284
rect 3265 264 3269 284
rect 3325 264 3329 304
rect 3345 264 3349 304
rect 3365 264 3369 304
rect 3432 264 3436 284
rect 3454 264 3458 304
rect 3462 264 3466 304
rect 3525 264 3529 284
rect 3545 264 3549 284
rect 3591 264 3595 284
rect 3611 264 3615 284
rect 3631 264 3635 304
rect 3693 264 3697 304
rect 3703 264 3707 304
rect 3773 264 3777 304
rect 3783 264 3787 304
rect 3865 264 3869 304
rect 3885 264 3889 304
rect 3905 264 3909 304
rect 3965 264 3969 284
rect 4025 264 4029 284
rect 4071 264 4075 304
rect 4093 264 4097 284
rect 4103 264 4107 284
rect 4123 264 4127 284
rect 4131 264 4135 284
rect 4177 264 4181 284
rect 4199 264 4203 284
rect 4209 264 4213 284
rect 4231 264 4235 284
rect 4241 264 4245 284
rect 4261 264 4265 304
rect 4333 264 4337 304
rect 4343 264 4347 304
rect 4405 264 4409 304
rect 4425 264 4429 304
rect 4445 264 4449 304
rect 4505 264 4509 284
rect 4551 264 4555 304
rect 4573 264 4577 284
rect 4583 264 4587 284
rect 4603 264 4607 284
rect 4611 264 4615 284
rect 4657 264 4661 284
rect 4679 264 4683 284
rect 4689 264 4693 284
rect 4711 264 4715 284
rect 4721 264 4725 284
rect 4741 264 4745 304
rect 68 176 72 236
rect 76 176 80 236
rect 84 176 88 236
rect 134 196 138 236
rect 142 196 146 236
rect 164 216 168 236
rect 245 196 249 236
rect 265 196 269 236
rect 285 196 289 236
rect 331 196 335 236
rect 351 196 355 236
rect 371 196 375 236
rect 468 176 472 236
rect 476 176 480 236
rect 484 176 488 236
rect 532 176 536 236
rect 540 176 544 236
rect 548 176 552 236
rect 634 196 638 236
rect 642 196 646 236
rect 664 216 668 236
rect 752 216 756 236
rect 774 196 778 236
rect 782 196 786 236
rect 831 216 835 236
rect 905 196 909 236
rect 925 196 929 236
rect 945 196 949 236
rect 1005 216 1009 236
rect 1051 196 1055 236
rect 1071 196 1075 236
rect 1091 196 1095 236
rect 1151 196 1155 236
rect 1171 196 1175 236
rect 1191 196 1195 236
rect 1252 176 1256 236
rect 1260 176 1264 236
rect 1268 176 1272 236
rect 1352 176 1356 236
rect 1360 176 1364 236
rect 1368 176 1372 236
rect 1472 216 1476 236
rect 1494 196 1498 236
rect 1502 196 1506 236
rect 1552 176 1556 236
rect 1560 176 1564 236
rect 1568 176 1572 236
rect 1672 216 1676 236
rect 1694 196 1698 236
rect 1702 196 1706 236
rect 1752 176 1756 236
rect 1760 176 1764 236
rect 1768 176 1772 236
rect 1853 196 1857 236
rect 1863 196 1867 236
rect 1931 216 1935 236
rect 1953 196 1957 236
rect 2035 196 2039 236
rect 2055 196 2059 236
rect 2065 196 2069 236
rect 2111 216 2115 236
rect 2133 196 2137 236
rect 2192 176 2196 236
rect 2200 176 2204 236
rect 2208 176 2212 236
rect 2294 196 2298 236
rect 2302 196 2306 236
rect 2322 196 2326 236
rect 2330 196 2334 236
rect 2411 196 2415 236
rect 2431 196 2435 236
rect 2451 196 2455 236
rect 2532 216 2536 236
rect 2554 196 2558 236
rect 2562 196 2566 236
rect 2611 196 2615 236
rect 2631 196 2635 236
rect 2651 196 2655 236
rect 2711 216 2715 236
rect 2772 176 2776 236
rect 2780 176 2784 236
rect 2788 176 2792 236
rect 2871 216 2875 236
rect 2935 196 2939 236
rect 2955 216 2959 236
rect 2965 216 2969 236
rect 2987 216 2991 236
rect 2997 216 3001 236
rect 3019 216 3023 236
rect 3065 216 3069 236
rect 3073 216 3077 236
rect 3093 216 3097 236
rect 3103 216 3107 236
rect 3125 196 3129 236
rect 3171 216 3175 236
rect 3245 216 3249 236
rect 3295 196 3299 236
rect 3315 216 3319 236
rect 3325 216 3329 236
rect 3347 216 3351 236
rect 3357 216 3361 236
rect 3379 216 3383 236
rect 3425 216 3429 236
rect 3433 216 3437 236
rect 3453 216 3457 236
rect 3463 216 3467 236
rect 3485 196 3489 236
rect 3545 216 3549 236
rect 3565 216 3569 236
rect 3611 196 3615 236
rect 3633 216 3637 236
rect 3643 216 3647 236
rect 3663 216 3667 236
rect 3671 216 3675 236
rect 3717 216 3721 236
rect 3739 216 3743 236
rect 3749 216 3753 236
rect 3771 216 3775 236
rect 3781 216 3785 236
rect 3801 196 3805 236
rect 3851 216 3855 236
rect 3911 196 3915 236
rect 3931 196 3935 236
rect 3951 196 3955 236
rect 4011 216 4015 236
rect 4031 216 4035 236
rect 4091 216 4095 236
rect 4111 216 4115 236
rect 4185 216 4189 236
rect 4205 216 4209 236
rect 4251 196 4255 236
rect 4271 196 4275 236
rect 4291 196 4295 236
rect 4373 196 4377 236
rect 4383 196 4387 236
rect 4445 216 4449 236
rect 4491 216 4495 236
rect 4511 216 4515 236
rect 4573 196 4577 236
rect 4583 196 4587 236
rect 4665 216 4669 236
rect 4713 196 4717 236
rect 4723 196 4727 236
<< ptransistor >>
rect 45 4344 49 4424
rect 65 4344 69 4424
rect 85 4344 89 4424
rect 145 4344 149 4384
rect 165 4344 169 4384
rect 185 4344 189 4384
rect 231 4344 235 4384
rect 251 4344 255 4384
rect 271 4344 275 4384
rect 345 4344 349 4384
rect 365 4344 369 4384
rect 385 4344 389 4384
rect 431 4344 435 4424
rect 451 4344 455 4424
rect 471 4344 475 4424
rect 536 4344 540 4424
rect 544 4344 548 4424
rect 566 4344 570 4384
rect 636 4344 640 4424
rect 644 4344 648 4424
rect 666 4344 670 4384
rect 745 4344 749 4384
rect 765 4344 769 4384
rect 785 4344 789 4384
rect 831 4344 835 4384
rect 851 4344 855 4384
rect 871 4344 875 4384
rect 931 4344 935 4384
rect 951 4344 955 4384
rect 1011 4344 1015 4384
rect 1031 4344 1035 4384
rect 1051 4344 1055 4384
rect 1111 4344 1115 4424
rect 1131 4344 1135 4424
rect 1151 4344 1155 4424
rect 1225 4344 1229 4384
rect 1245 4344 1249 4384
rect 1317 4344 1321 4424
rect 1325 4344 1329 4424
rect 1390 4344 1394 4384
rect 1412 4344 1416 4424
rect 1420 4344 1424 4424
rect 1485 4344 1489 4384
rect 1505 4344 1509 4384
rect 1551 4344 1555 4424
rect 1559 4344 1563 4424
rect 1631 4344 1635 4384
rect 1651 4344 1655 4384
rect 1671 4344 1675 4384
rect 1745 4344 1749 4424
rect 1765 4344 1769 4424
rect 1785 4344 1789 4424
rect 1831 4344 1835 4384
rect 1905 4344 1909 4384
rect 1951 4344 1955 4424
rect 1971 4344 1975 4424
rect 1991 4344 1995 4424
rect 2051 4344 2055 4424
rect 2059 4344 2063 4424
rect 2131 4344 2135 4384
rect 2196 4344 2200 4424
rect 2204 4344 2208 4424
rect 2226 4344 2230 4384
rect 2315 4344 2319 4424
rect 2325 4344 2329 4424
rect 2355 4344 2359 4424
rect 2365 4344 2369 4424
rect 2411 4344 2415 4424
rect 2421 4344 2425 4424
rect 2441 4344 2445 4424
rect 2511 4344 2515 4424
rect 2531 4344 2535 4424
rect 2551 4344 2555 4424
rect 2625 4344 2629 4424
rect 2645 4344 2649 4424
rect 2665 4344 2669 4424
rect 2685 4344 2689 4424
rect 2735 4344 2739 4424
rect 2755 4344 2759 4384
rect 2769 4344 2773 4384
rect 2789 4344 2793 4384
rect 2801 4344 2805 4384
rect 2821 4344 2825 4384
rect 2867 4344 2871 4384
rect 2875 4344 2879 4384
rect 2895 4344 2899 4364
rect 2903 4344 2907 4364
rect 2925 4344 2929 4424
rect 2985 4344 2989 4384
rect 3050 4344 3054 4384
rect 3072 4344 3076 4424
rect 3080 4344 3084 4424
rect 3157 4344 3161 4424
rect 3165 4344 3169 4424
rect 3230 4344 3234 4384
rect 3252 4344 3256 4424
rect 3260 4344 3264 4424
rect 3337 4344 3341 4424
rect 3345 4344 3349 4424
rect 3405 4344 3409 4384
rect 3451 4344 3455 4424
rect 3473 4344 3477 4364
rect 3481 4344 3485 4364
rect 3501 4344 3505 4384
rect 3509 4344 3513 4384
rect 3555 4344 3559 4384
rect 3575 4344 3579 4384
rect 3587 4344 3591 4384
rect 3607 4344 3611 4384
rect 3621 4344 3625 4384
rect 3641 4344 3645 4424
rect 3696 4344 3700 4424
rect 3704 4344 3708 4424
rect 3726 4344 3730 4384
rect 3791 4344 3795 4384
rect 3811 4344 3815 4384
rect 3885 4344 3889 4424
rect 3905 4344 3909 4424
rect 3925 4344 3929 4424
rect 3945 4344 3949 4424
rect 3965 4344 3969 4424
rect 3985 4344 3989 4424
rect 4005 4344 4009 4424
rect 4025 4344 4029 4424
rect 4083 4344 4087 4424
rect 4105 4344 4109 4384
rect 4151 4344 4155 4384
rect 4171 4344 4175 4384
rect 4231 4344 4235 4384
rect 4296 4344 4300 4424
rect 4304 4344 4308 4424
rect 4326 4344 4330 4384
rect 4391 4344 4395 4424
rect 4413 4344 4417 4364
rect 4421 4344 4425 4364
rect 4441 4344 4445 4384
rect 4449 4344 4453 4384
rect 4495 4344 4499 4384
rect 4515 4344 4519 4384
rect 4527 4344 4531 4384
rect 4547 4344 4551 4384
rect 4561 4344 4565 4384
rect 4581 4344 4585 4424
rect 4631 4344 4635 4384
rect 4653 4344 4657 4424
rect 4711 4344 4715 4384
rect 4731 4344 4735 4384
rect 45 4276 49 4316
rect 65 4276 69 4316
rect 111 4236 115 4316
rect 131 4236 135 4316
rect 151 4236 155 4316
rect 225 4276 229 4316
rect 245 4276 249 4316
rect 317 4236 321 4316
rect 325 4236 329 4316
rect 390 4276 394 4316
rect 412 4236 416 4316
rect 420 4236 424 4316
rect 476 4236 480 4316
rect 484 4236 488 4316
rect 506 4276 510 4316
rect 585 4276 589 4316
rect 645 4236 649 4316
rect 665 4236 669 4316
rect 685 4236 689 4316
rect 745 4276 749 4316
rect 791 4276 795 4316
rect 811 4276 815 4316
rect 831 4276 835 4316
rect 905 4236 909 4316
rect 925 4236 929 4316
rect 945 4236 949 4316
rect 965 4236 969 4316
rect 1025 4276 1029 4316
rect 1045 4276 1049 4316
rect 1065 4276 1069 4316
rect 1111 4276 1115 4316
rect 1131 4276 1135 4316
rect 1151 4276 1155 4316
rect 1225 4276 1229 4316
rect 1245 4276 1249 4316
rect 1305 4276 1309 4316
rect 1325 4276 1329 4316
rect 1345 4276 1349 4316
rect 1405 4276 1409 4316
rect 1425 4276 1429 4316
rect 1471 4276 1475 4316
rect 1491 4276 1495 4316
rect 1511 4276 1515 4316
rect 1597 4236 1601 4316
rect 1605 4236 1609 4316
rect 1677 4236 1681 4316
rect 1685 4236 1689 4316
rect 1736 4236 1740 4316
rect 1744 4236 1748 4316
rect 1766 4276 1770 4316
rect 1845 4276 1849 4316
rect 1865 4276 1869 4316
rect 1911 4276 1915 4316
rect 1971 4276 1975 4316
rect 1991 4276 1995 4316
rect 2011 4276 2015 4316
rect 2071 4276 2075 4316
rect 2091 4276 2095 4316
rect 2111 4276 2115 4316
rect 2175 4236 2179 4316
rect 2195 4276 2199 4316
rect 2209 4276 2213 4316
rect 2229 4276 2233 4316
rect 2241 4276 2245 4316
rect 2261 4276 2265 4316
rect 2307 4276 2311 4316
rect 2315 4276 2319 4316
rect 2335 4296 2339 4316
rect 2343 4296 2347 4316
rect 2365 4236 2369 4316
rect 2411 4276 2415 4316
rect 2433 4236 2437 4316
rect 2505 4276 2509 4316
rect 2577 4236 2581 4316
rect 2585 4236 2589 4316
rect 2631 4236 2635 4316
rect 2653 4296 2657 4316
rect 2661 4296 2665 4316
rect 2681 4276 2685 4316
rect 2689 4276 2693 4316
rect 2735 4276 2739 4316
rect 2755 4276 2759 4316
rect 2767 4276 2771 4316
rect 2787 4276 2791 4316
rect 2801 4276 2805 4316
rect 2821 4236 2825 4316
rect 2871 4276 2875 4316
rect 2957 4236 2961 4316
rect 2965 4236 2969 4316
rect 3016 4236 3020 4316
rect 3024 4236 3028 4316
rect 3046 4276 3050 4316
rect 3111 4276 3115 4316
rect 3131 4276 3135 4316
rect 3205 4276 3209 4316
rect 3225 4276 3229 4316
rect 3285 4276 3289 4316
rect 3305 4276 3309 4316
rect 3351 4236 3355 4316
rect 3359 4236 3363 4316
rect 3435 4236 3439 4316
rect 3455 4276 3459 4316
rect 3469 4276 3473 4316
rect 3489 4276 3493 4316
rect 3501 4276 3505 4316
rect 3521 4276 3525 4316
rect 3567 4276 3571 4316
rect 3575 4276 3579 4316
rect 3595 4296 3599 4316
rect 3603 4296 3607 4316
rect 3625 4236 3629 4316
rect 3685 4276 3689 4316
rect 3705 4276 3709 4316
rect 3751 4236 3755 4316
rect 3759 4236 3763 4316
rect 3831 4236 3835 4316
rect 3853 4296 3857 4316
rect 3861 4296 3865 4316
rect 3881 4276 3885 4316
rect 3889 4276 3893 4316
rect 3935 4276 3939 4316
rect 3955 4276 3959 4316
rect 3967 4276 3971 4316
rect 3987 4276 3991 4316
rect 4001 4276 4005 4316
rect 4021 4236 4025 4316
rect 4071 4236 4075 4316
rect 4079 4236 4083 4316
rect 4165 4236 4169 4316
rect 4185 4236 4189 4316
rect 4205 4236 4209 4316
rect 4251 4276 4255 4316
rect 4273 4236 4277 4316
rect 4357 4236 4361 4316
rect 4365 4236 4369 4316
rect 4425 4236 4429 4316
rect 4445 4236 4449 4316
rect 4465 4236 4469 4316
rect 4511 4236 4515 4316
rect 4533 4296 4537 4316
rect 4541 4296 4545 4316
rect 4561 4276 4565 4316
rect 4569 4276 4573 4316
rect 4615 4276 4619 4316
rect 4635 4276 4639 4316
rect 4647 4276 4651 4316
rect 4667 4276 4671 4316
rect 4681 4276 4685 4316
rect 4701 4236 4705 4316
rect 45 3864 49 3904
rect 65 3864 69 3904
rect 111 3864 115 3904
rect 131 3864 135 3904
rect 205 3864 209 3904
rect 225 3864 229 3904
rect 290 3864 294 3904
rect 312 3864 316 3944
rect 320 3864 324 3944
rect 371 3864 375 3944
rect 391 3864 395 3944
rect 411 3864 415 3944
rect 497 3864 501 3944
rect 505 3864 509 3944
rect 551 3864 555 3904
rect 571 3864 575 3904
rect 636 3864 640 3944
rect 644 3864 648 3944
rect 666 3864 670 3904
rect 745 3864 749 3904
rect 765 3864 769 3904
rect 785 3864 789 3904
rect 831 3864 835 3904
rect 851 3864 855 3904
rect 871 3864 875 3904
rect 950 3864 954 3904
rect 972 3864 976 3944
rect 980 3864 984 3944
rect 1036 3864 1040 3944
rect 1044 3864 1048 3944
rect 1066 3864 1070 3904
rect 1145 3864 1149 3904
rect 1205 3864 1209 3904
rect 1225 3864 1229 3904
rect 1245 3864 1249 3904
rect 1291 3864 1295 3904
rect 1351 3864 1355 3904
rect 1371 3864 1375 3904
rect 1391 3864 1395 3904
rect 1451 3864 1455 3904
rect 1471 3864 1475 3904
rect 1491 3864 1495 3904
rect 1551 3864 1555 3904
rect 1571 3864 1575 3904
rect 1657 3864 1661 3944
rect 1665 3864 1669 3944
rect 1721 3864 1725 3944
rect 1743 3864 1747 3904
rect 1765 3864 1769 3904
rect 1830 3864 1834 3904
rect 1852 3864 1856 3944
rect 1860 3864 1864 3944
rect 1911 3864 1915 3944
rect 1919 3864 1923 3944
rect 2005 3864 2009 3904
rect 2056 3864 2060 3944
rect 2064 3864 2068 3944
rect 2086 3864 2090 3904
rect 2151 3864 2155 3904
rect 2211 3864 2215 3904
rect 2231 3864 2235 3904
rect 2291 3864 2295 3904
rect 2311 3864 2315 3904
rect 2331 3864 2335 3904
rect 2391 3864 2395 3904
rect 2413 3864 2417 3944
rect 2471 3864 2475 3944
rect 2491 3864 2495 3944
rect 2511 3864 2515 3944
rect 2531 3864 2535 3944
rect 2551 3864 2555 3944
rect 2571 3864 2575 3944
rect 2591 3864 2595 3944
rect 2611 3864 2615 3944
rect 2675 3864 2679 3944
rect 2695 3864 2699 3904
rect 2709 3864 2713 3904
rect 2729 3864 2733 3904
rect 2741 3864 2745 3904
rect 2761 3864 2765 3904
rect 2807 3864 2811 3904
rect 2815 3864 2819 3904
rect 2835 3864 2839 3884
rect 2843 3864 2847 3884
rect 2865 3864 2869 3944
rect 2911 3864 2915 3904
rect 2976 3864 2980 3944
rect 2984 3864 2988 3944
rect 3006 3864 3010 3904
rect 3071 3864 3075 3944
rect 3079 3864 3083 3944
rect 3151 3864 3155 3904
rect 3171 3864 3175 3904
rect 3245 3864 3249 3944
rect 3265 3864 3269 3944
rect 3285 3864 3289 3944
rect 3331 3864 3335 3904
rect 3353 3864 3357 3904
rect 3375 3864 3379 3944
rect 3457 3864 3461 3944
rect 3465 3864 3469 3944
rect 3525 3864 3529 3904
rect 3571 3864 3575 3944
rect 3593 3864 3597 3884
rect 3601 3864 3605 3884
rect 3621 3864 3625 3904
rect 3629 3864 3633 3904
rect 3675 3864 3679 3904
rect 3695 3864 3699 3904
rect 3707 3864 3711 3904
rect 3727 3864 3731 3904
rect 3741 3864 3745 3904
rect 3761 3864 3765 3944
rect 3825 3864 3829 3944
rect 3845 3864 3849 3944
rect 3865 3864 3869 3944
rect 3911 3864 3915 3944
rect 3919 3864 3923 3944
rect 4017 3864 4021 3944
rect 4025 3864 4029 3944
rect 4071 3864 4075 3904
rect 4093 3864 4097 3904
rect 4115 3864 4119 3944
rect 4176 3864 4180 3944
rect 4184 3864 4188 3944
rect 4206 3864 4210 3904
rect 4290 3864 4294 3904
rect 4312 3864 4316 3944
rect 4320 3864 4324 3944
rect 4385 3864 4389 3904
rect 4431 3864 4435 3944
rect 4453 3864 4457 3884
rect 4461 3864 4465 3884
rect 4481 3864 4485 3904
rect 4489 3864 4493 3904
rect 4535 3864 4539 3904
rect 4555 3864 4559 3904
rect 4567 3864 4571 3904
rect 4587 3864 4591 3904
rect 4601 3864 4605 3904
rect 4621 3864 4625 3944
rect 4671 3864 4675 3904
rect 57 3756 61 3836
rect 65 3756 69 3836
rect 116 3756 120 3836
rect 124 3756 128 3836
rect 146 3796 150 3836
rect 225 3796 229 3836
rect 285 3756 289 3836
rect 305 3756 309 3836
rect 325 3756 329 3836
rect 381 3756 385 3836
rect 403 3796 407 3836
rect 425 3796 429 3836
rect 485 3796 489 3836
rect 505 3796 509 3836
rect 565 3796 569 3836
rect 585 3796 589 3836
rect 631 3796 635 3836
rect 696 3756 700 3836
rect 704 3756 708 3836
rect 726 3796 730 3836
rect 791 3796 795 3836
rect 811 3796 815 3836
rect 885 3796 889 3836
rect 905 3796 909 3836
rect 925 3796 929 3836
rect 971 3756 975 3836
rect 991 3756 995 3836
rect 1011 3756 1015 3836
rect 1071 3796 1075 3836
rect 1091 3796 1095 3836
rect 1111 3796 1115 3836
rect 1171 3756 1175 3836
rect 1191 3756 1195 3836
rect 1211 3756 1215 3836
rect 1271 3796 1275 3836
rect 1345 3796 1349 3836
rect 1365 3796 1369 3836
rect 1385 3796 1389 3836
rect 1445 3796 1449 3836
rect 1510 3796 1514 3836
rect 1532 3756 1536 3836
rect 1540 3756 1544 3836
rect 1605 3796 1609 3836
rect 1651 3756 1655 3836
rect 1671 3756 1675 3836
rect 1691 3756 1695 3836
rect 1751 3756 1755 3836
rect 1759 3756 1763 3836
rect 1845 3756 1849 3836
rect 1865 3756 1869 3836
rect 1885 3756 1889 3836
rect 1945 3796 1949 3836
rect 1965 3796 1969 3836
rect 2011 3756 2015 3836
rect 2021 3756 2025 3836
rect 2041 3756 2045 3836
rect 2111 3796 2115 3836
rect 2133 3756 2137 3836
rect 2205 3756 2209 3836
rect 2225 3756 2229 3836
rect 2245 3756 2249 3836
rect 2265 3756 2269 3836
rect 2285 3756 2289 3836
rect 2305 3756 2309 3836
rect 2325 3756 2329 3836
rect 2345 3756 2349 3836
rect 2395 3756 2399 3836
rect 2415 3796 2419 3836
rect 2429 3796 2433 3836
rect 2449 3796 2453 3836
rect 2461 3796 2465 3836
rect 2481 3796 2485 3836
rect 2527 3796 2531 3836
rect 2535 3796 2539 3836
rect 2555 3816 2559 3836
rect 2563 3816 2567 3836
rect 2585 3756 2589 3836
rect 2650 3796 2654 3836
rect 2672 3756 2676 3836
rect 2680 3756 2684 3836
rect 2745 3796 2749 3836
rect 2817 3756 2821 3836
rect 2825 3756 2829 3836
rect 2897 3756 2901 3836
rect 2905 3756 2909 3836
rect 2977 3756 2981 3836
rect 2985 3756 2989 3836
rect 3031 3796 3035 3836
rect 3105 3796 3109 3836
rect 3156 3756 3160 3836
rect 3164 3756 3168 3836
rect 3186 3796 3190 3836
rect 3265 3756 3269 3836
rect 3285 3756 3289 3836
rect 3305 3756 3309 3836
rect 3351 3756 3355 3836
rect 3371 3756 3375 3836
rect 3391 3756 3395 3836
rect 3451 3796 3455 3836
rect 3511 3796 3515 3836
rect 3533 3796 3537 3836
rect 3555 3756 3559 3836
rect 3616 3756 3620 3836
rect 3624 3756 3628 3836
rect 3646 3796 3650 3836
rect 3716 3756 3720 3836
rect 3724 3756 3728 3836
rect 3746 3796 3750 3836
rect 3815 3756 3819 3836
rect 3835 3796 3839 3836
rect 3849 3796 3853 3836
rect 3869 3796 3873 3836
rect 3881 3796 3885 3836
rect 3901 3796 3905 3836
rect 3947 3796 3951 3836
rect 3955 3796 3959 3836
rect 3975 3816 3979 3836
rect 3983 3816 3987 3836
rect 4005 3756 4009 3836
rect 4051 3796 4055 3836
rect 4073 3756 4077 3836
rect 4157 3756 4161 3836
rect 4165 3756 4169 3836
rect 4211 3756 4215 3836
rect 4231 3756 4235 3836
rect 4251 3756 4255 3836
rect 4311 3756 4315 3836
rect 4333 3816 4337 3836
rect 4341 3816 4345 3836
rect 4361 3796 4365 3836
rect 4369 3796 4373 3836
rect 4415 3796 4419 3836
rect 4435 3796 4439 3836
rect 4447 3796 4451 3836
rect 4467 3796 4471 3836
rect 4481 3796 4485 3836
rect 4501 3756 4505 3836
rect 4551 3796 4555 3836
rect 4573 3756 4577 3836
rect 4645 3796 4649 3836
rect 4691 3796 4695 3836
rect 45 3384 49 3424
rect 65 3384 69 3424
rect 115 3384 119 3464
rect 135 3384 139 3424
rect 149 3384 153 3424
rect 169 3384 173 3424
rect 181 3384 185 3424
rect 201 3384 205 3424
rect 247 3384 251 3424
rect 255 3384 259 3424
rect 275 3384 279 3404
rect 283 3384 287 3404
rect 305 3384 309 3464
rect 365 3384 369 3424
rect 425 3384 429 3424
rect 445 3384 449 3424
rect 510 3384 514 3424
rect 532 3384 536 3464
rect 540 3384 544 3464
rect 610 3384 614 3424
rect 632 3384 636 3464
rect 640 3384 644 3464
rect 691 3384 695 3424
rect 711 3384 715 3424
rect 771 3384 775 3464
rect 781 3384 785 3464
rect 811 3384 815 3464
rect 821 3384 825 3464
rect 891 3384 895 3424
rect 965 3384 969 3424
rect 985 3384 989 3424
rect 1005 3384 1009 3424
rect 1051 3384 1055 3464
rect 1071 3384 1075 3464
rect 1091 3384 1095 3464
rect 1151 3384 1155 3464
rect 1159 3384 1163 3464
rect 1231 3384 1235 3424
rect 1251 3384 1255 3424
rect 1311 3384 1315 3424
rect 1331 3384 1335 3424
rect 1396 3384 1400 3464
rect 1404 3384 1408 3464
rect 1426 3384 1430 3424
rect 1495 3384 1499 3464
rect 1515 3384 1519 3424
rect 1529 3384 1533 3424
rect 1549 3384 1553 3424
rect 1561 3384 1565 3424
rect 1581 3384 1585 3424
rect 1627 3384 1631 3424
rect 1635 3384 1639 3424
rect 1655 3384 1659 3404
rect 1663 3384 1667 3404
rect 1685 3384 1689 3464
rect 1745 3384 1749 3424
rect 1765 3384 1769 3424
rect 1816 3384 1820 3464
rect 1824 3384 1828 3464
rect 1846 3384 1850 3424
rect 1911 3384 1915 3464
rect 1985 3384 1989 3424
rect 2005 3384 2009 3424
rect 2061 3384 2065 3464
rect 2083 3384 2087 3424
rect 2105 3384 2109 3424
rect 2151 3384 2155 3424
rect 2171 3384 2175 3424
rect 2231 3384 2235 3424
rect 2251 3384 2255 3424
rect 2271 3384 2275 3424
rect 2331 3384 2335 3424
rect 2391 3384 2395 3424
rect 2451 3384 2455 3464
rect 2473 3384 2477 3404
rect 2481 3384 2485 3404
rect 2501 3384 2505 3424
rect 2509 3384 2513 3424
rect 2555 3384 2559 3424
rect 2575 3384 2579 3424
rect 2587 3384 2591 3424
rect 2607 3384 2611 3424
rect 2621 3384 2625 3424
rect 2641 3384 2645 3464
rect 2696 3384 2700 3464
rect 2704 3384 2708 3464
rect 2726 3384 2730 3424
rect 2791 3384 2795 3424
rect 2813 3384 2817 3464
rect 2871 3384 2875 3424
rect 2891 3384 2895 3424
rect 2951 3384 2955 3464
rect 2973 3384 2977 3404
rect 2981 3384 2985 3404
rect 3001 3384 3005 3424
rect 3009 3384 3013 3424
rect 3055 3384 3059 3424
rect 3075 3384 3079 3424
rect 3087 3384 3091 3424
rect 3107 3384 3111 3424
rect 3121 3384 3125 3424
rect 3141 3384 3145 3464
rect 3210 3384 3214 3424
rect 3232 3384 3236 3464
rect 3240 3384 3244 3464
rect 3305 3384 3309 3424
rect 3351 3384 3355 3464
rect 3359 3384 3363 3464
rect 3431 3384 3435 3424
rect 3517 3384 3521 3464
rect 3525 3384 3529 3464
rect 3571 3384 3575 3464
rect 3591 3384 3595 3464
rect 3611 3384 3615 3464
rect 3671 3384 3675 3464
rect 3681 3384 3685 3464
rect 3701 3384 3705 3464
rect 3785 3384 3789 3464
rect 3805 3384 3809 3464
rect 3825 3384 3829 3464
rect 3845 3384 3849 3464
rect 3905 3384 3909 3424
rect 3925 3384 3929 3424
rect 3971 3384 3975 3464
rect 3993 3384 3997 3404
rect 4001 3384 4005 3404
rect 4021 3384 4025 3424
rect 4029 3384 4033 3424
rect 4075 3384 4079 3424
rect 4095 3384 4099 3424
rect 4107 3384 4111 3424
rect 4127 3384 4131 3424
rect 4141 3384 4145 3424
rect 4161 3384 4165 3464
rect 4211 3384 4215 3464
rect 4233 3384 4237 3404
rect 4241 3384 4245 3404
rect 4261 3384 4265 3424
rect 4269 3384 4273 3424
rect 4315 3384 4319 3424
rect 4335 3384 4339 3424
rect 4347 3384 4351 3424
rect 4367 3384 4371 3424
rect 4381 3384 4385 3424
rect 4401 3384 4405 3464
rect 4465 3384 4469 3464
rect 4485 3384 4489 3464
rect 4505 3384 4509 3464
rect 4525 3384 4529 3464
rect 4545 3384 4549 3464
rect 4565 3384 4569 3464
rect 4585 3384 4589 3464
rect 4605 3384 4609 3464
rect 4656 3384 4660 3464
rect 4664 3384 4668 3464
rect 4686 3384 4690 3424
rect 35 3276 39 3356
rect 55 3316 59 3356
rect 69 3316 73 3356
rect 89 3316 93 3356
rect 101 3316 105 3356
rect 121 3316 125 3356
rect 167 3316 171 3356
rect 175 3316 179 3356
rect 195 3336 199 3356
rect 203 3336 207 3356
rect 225 3276 229 3356
rect 285 3276 289 3356
rect 305 3276 309 3356
rect 325 3276 329 3356
rect 345 3276 349 3356
rect 405 3316 409 3356
rect 425 3316 429 3356
rect 471 3276 475 3356
rect 493 3336 497 3356
rect 501 3336 505 3356
rect 521 3316 525 3356
rect 529 3316 533 3356
rect 575 3316 579 3356
rect 595 3316 599 3356
rect 607 3316 611 3356
rect 627 3316 631 3356
rect 641 3316 645 3356
rect 661 3276 665 3356
rect 730 3316 734 3356
rect 752 3276 756 3356
rect 760 3276 764 3356
rect 825 3276 829 3356
rect 845 3276 849 3356
rect 865 3276 869 3356
rect 885 3276 889 3356
rect 931 3316 935 3356
rect 951 3316 955 3356
rect 1025 3316 1029 3356
rect 1045 3316 1049 3356
rect 1065 3316 1069 3356
rect 1121 3276 1125 3356
rect 1143 3316 1147 3356
rect 1165 3316 1169 3356
rect 1211 3316 1215 3356
rect 1231 3316 1235 3356
rect 1251 3316 1255 3356
rect 1316 3276 1320 3356
rect 1324 3276 1328 3356
rect 1346 3316 1350 3356
rect 1411 3316 1415 3356
rect 1431 3316 1435 3356
rect 1515 3276 1519 3356
rect 1535 3276 1539 3356
rect 1545 3276 1549 3356
rect 1605 3316 1609 3356
rect 1625 3316 1629 3356
rect 1676 3276 1680 3356
rect 1684 3276 1688 3356
rect 1706 3316 1710 3356
rect 1790 3316 1794 3356
rect 1812 3276 1816 3356
rect 1820 3276 1824 3356
rect 1871 3316 1875 3356
rect 1891 3316 1895 3356
rect 1956 3276 1960 3356
rect 1964 3276 1968 3356
rect 1986 3316 1990 3356
rect 2070 3316 2074 3356
rect 2092 3276 2096 3356
rect 2100 3276 2104 3356
rect 2151 3316 2155 3356
rect 2216 3276 2220 3356
rect 2224 3276 2228 3356
rect 2246 3316 2250 3356
rect 2325 3316 2329 3356
rect 2371 3316 2375 3356
rect 2391 3316 2395 3356
rect 2451 3276 2455 3356
rect 2473 3336 2477 3356
rect 2481 3336 2485 3356
rect 2501 3316 2505 3356
rect 2509 3316 2513 3356
rect 2555 3316 2559 3356
rect 2575 3316 2579 3356
rect 2587 3316 2591 3356
rect 2607 3316 2611 3356
rect 2621 3316 2625 3356
rect 2641 3276 2645 3356
rect 2691 3316 2695 3356
rect 2713 3276 2717 3356
rect 2771 3276 2775 3356
rect 2793 3336 2797 3356
rect 2801 3336 2805 3356
rect 2821 3316 2825 3356
rect 2829 3316 2833 3356
rect 2875 3316 2879 3356
rect 2895 3316 2899 3356
rect 2907 3316 2911 3356
rect 2927 3316 2931 3356
rect 2941 3316 2945 3356
rect 2961 3276 2965 3356
rect 3030 3316 3034 3356
rect 3052 3276 3056 3356
rect 3060 3276 3064 3356
rect 3130 3316 3134 3356
rect 3152 3276 3156 3356
rect 3160 3276 3164 3356
rect 3216 3276 3220 3356
rect 3224 3276 3228 3356
rect 3246 3316 3250 3356
rect 3330 3316 3334 3356
rect 3352 3276 3356 3356
rect 3360 3276 3364 3356
rect 3416 3276 3420 3356
rect 3424 3276 3428 3356
rect 3446 3316 3450 3356
rect 3511 3316 3515 3356
rect 3531 3316 3535 3356
rect 3591 3316 3595 3356
rect 3611 3316 3615 3356
rect 3671 3316 3675 3356
rect 3691 3316 3695 3356
rect 3751 3316 3755 3356
rect 3771 3316 3775 3356
rect 3831 3316 3835 3356
rect 3853 3276 3857 3356
rect 3925 3316 3929 3356
rect 3945 3316 3949 3356
rect 4017 3276 4021 3356
rect 4025 3276 4029 3356
rect 4071 3316 4075 3356
rect 4093 3276 4097 3356
rect 4165 3316 4169 3356
rect 4230 3316 4234 3356
rect 4252 3276 4256 3356
rect 4260 3276 4264 3356
rect 4325 3316 4329 3356
rect 4376 3276 4380 3356
rect 4384 3276 4388 3356
rect 4406 3316 4410 3356
rect 4485 3316 4489 3356
rect 4505 3316 4509 3356
rect 4555 3276 4559 3356
rect 4575 3316 4579 3356
rect 4589 3316 4593 3356
rect 4609 3316 4613 3356
rect 4621 3316 4625 3356
rect 4641 3316 4645 3356
rect 4687 3316 4691 3356
rect 4695 3316 4699 3356
rect 4715 3336 4719 3356
rect 4723 3336 4727 3356
rect 4745 3276 4749 3356
rect 45 2904 49 2984
rect 65 2904 69 2984
rect 85 2904 89 2984
rect 105 2904 109 2984
rect 161 2904 165 2984
rect 183 2904 187 2944
rect 205 2904 209 2944
rect 251 2904 255 2984
rect 273 2904 277 2924
rect 281 2904 285 2924
rect 301 2904 305 2944
rect 309 2904 313 2944
rect 355 2904 359 2944
rect 375 2904 379 2944
rect 387 2904 391 2944
rect 407 2904 411 2944
rect 421 2904 425 2944
rect 441 2904 445 2984
rect 496 2904 500 2984
rect 504 2904 508 2984
rect 526 2904 530 2944
rect 591 2904 595 2944
rect 611 2904 615 2944
rect 685 2904 689 2944
rect 705 2904 709 2944
rect 777 2904 781 2984
rect 785 2904 789 2984
rect 831 2904 835 2944
rect 851 2904 855 2944
rect 930 2904 934 2944
rect 952 2904 956 2984
rect 960 2904 964 2984
rect 1030 2904 1034 2944
rect 1052 2904 1056 2984
rect 1060 2904 1064 2984
rect 1137 2904 1141 2984
rect 1145 2904 1149 2984
rect 1210 2904 1214 2944
rect 1232 2904 1236 2984
rect 1240 2904 1244 2984
rect 1291 2904 1295 2944
rect 1311 2904 1315 2944
rect 1385 2904 1389 2984
rect 1431 2904 1435 2944
rect 1451 2904 1455 2944
rect 1511 2904 1515 2944
rect 1531 2904 1535 2944
rect 1591 2904 1595 2944
rect 1613 2904 1617 2984
rect 1676 2904 1680 2984
rect 1684 2904 1688 2984
rect 1706 2904 1710 2944
rect 1776 2904 1780 2984
rect 1784 2904 1788 2984
rect 1806 2904 1810 2944
rect 1871 2904 1875 2984
rect 1879 2904 1883 2984
rect 1951 2904 1955 2984
rect 1971 2904 1975 2984
rect 1991 2904 1995 2984
rect 2051 2904 2055 2944
rect 2116 2904 2120 2984
rect 2124 2904 2128 2984
rect 2146 2904 2150 2944
rect 2211 2904 2215 2984
rect 2219 2904 2223 2984
rect 2305 2904 2309 2944
rect 2325 2904 2329 2944
rect 2376 2904 2380 2984
rect 2384 2904 2388 2984
rect 2406 2904 2410 2944
rect 2471 2904 2475 2944
rect 2536 2904 2540 2984
rect 2544 2904 2548 2984
rect 2566 2904 2570 2944
rect 2631 2904 2635 2944
rect 2653 2904 2657 2984
rect 2711 2904 2715 2944
rect 2731 2904 2735 2944
rect 2795 2904 2799 2984
rect 2815 2904 2819 2944
rect 2829 2904 2833 2944
rect 2849 2904 2853 2944
rect 2861 2904 2865 2944
rect 2881 2904 2885 2944
rect 2927 2904 2931 2944
rect 2935 2904 2939 2944
rect 2955 2904 2959 2924
rect 2963 2904 2967 2924
rect 2985 2904 2989 2984
rect 3057 2904 3061 2984
rect 3065 2904 3069 2984
rect 3125 2904 3129 2984
rect 3145 2904 3149 2984
rect 3165 2904 3169 2984
rect 3211 2904 3215 2984
rect 3219 2904 3223 2984
rect 3295 2904 3299 2984
rect 3315 2904 3319 2944
rect 3329 2904 3333 2944
rect 3349 2904 3353 2944
rect 3361 2904 3365 2944
rect 3381 2904 3385 2944
rect 3427 2904 3431 2944
rect 3435 2904 3439 2944
rect 3455 2904 3459 2924
rect 3463 2904 3467 2924
rect 3485 2904 3489 2984
rect 3535 2904 3539 2984
rect 3555 2904 3559 2944
rect 3569 2904 3573 2944
rect 3589 2904 3593 2944
rect 3601 2904 3605 2944
rect 3621 2904 3625 2944
rect 3667 2904 3671 2944
rect 3675 2904 3679 2944
rect 3695 2904 3699 2924
rect 3703 2904 3707 2924
rect 3725 2904 3729 2984
rect 3771 2904 3775 2984
rect 3779 2904 3783 2984
rect 3870 2904 3874 2944
rect 3892 2904 3896 2984
rect 3900 2904 3904 2984
rect 3970 2904 3974 2944
rect 3992 2904 3996 2984
rect 4000 2904 4004 2984
rect 4056 2904 4060 2984
rect 4064 2904 4068 2984
rect 4086 2904 4090 2944
rect 4156 2904 4160 2984
rect 4164 2904 4168 2984
rect 4186 2904 4190 2944
rect 4251 2904 4255 2944
rect 4311 2904 4315 2944
rect 4331 2904 4335 2944
rect 4351 2904 4355 2944
rect 4411 2904 4415 2984
rect 4433 2904 4437 2924
rect 4441 2904 4445 2924
rect 4461 2904 4465 2944
rect 4469 2904 4473 2944
rect 4515 2904 4519 2944
rect 4535 2904 4539 2944
rect 4547 2904 4551 2944
rect 4567 2904 4571 2944
rect 4581 2904 4585 2944
rect 4601 2904 4605 2984
rect 4656 2904 4660 2984
rect 4664 2904 4668 2984
rect 4686 2904 4690 2944
rect 45 2836 49 2876
rect 110 2836 114 2876
rect 132 2796 136 2876
rect 140 2796 144 2876
rect 191 2796 195 2876
rect 211 2796 215 2876
rect 231 2796 235 2876
rect 251 2796 255 2876
rect 311 2836 315 2876
rect 331 2836 335 2876
rect 391 2836 395 2876
rect 413 2836 417 2876
rect 435 2796 439 2876
rect 510 2836 514 2876
rect 532 2796 536 2876
rect 540 2796 544 2876
rect 591 2836 595 2876
rect 611 2836 615 2876
rect 685 2796 689 2876
rect 745 2796 749 2876
rect 791 2836 795 2876
rect 811 2836 815 2876
rect 871 2836 875 2876
rect 893 2836 897 2876
rect 915 2796 919 2876
rect 990 2836 994 2876
rect 1012 2796 1016 2876
rect 1020 2796 1024 2876
rect 1071 2836 1075 2876
rect 1091 2836 1095 2876
rect 1170 2836 1174 2876
rect 1192 2796 1196 2876
rect 1200 2796 1204 2876
rect 1251 2796 1255 2876
rect 1273 2856 1277 2876
rect 1281 2856 1285 2876
rect 1301 2836 1305 2876
rect 1309 2836 1313 2876
rect 1355 2836 1359 2876
rect 1375 2836 1379 2876
rect 1387 2836 1391 2876
rect 1407 2836 1411 2876
rect 1421 2836 1425 2876
rect 1441 2796 1445 2876
rect 1503 2796 1507 2876
rect 1525 2836 1529 2876
rect 1575 2796 1579 2876
rect 1595 2836 1599 2876
rect 1609 2836 1613 2876
rect 1629 2836 1633 2876
rect 1641 2836 1645 2876
rect 1661 2836 1665 2876
rect 1707 2836 1711 2876
rect 1715 2836 1719 2876
rect 1735 2856 1739 2876
rect 1743 2856 1747 2876
rect 1765 2796 1769 2876
rect 1816 2796 1820 2876
rect 1824 2796 1828 2876
rect 1846 2836 1850 2876
rect 1911 2836 1915 2876
rect 1971 2796 1975 2876
rect 1981 2796 1985 2876
rect 2011 2796 2015 2876
rect 2021 2796 2025 2876
rect 2117 2796 2121 2876
rect 2125 2796 2129 2876
rect 2197 2796 2201 2876
rect 2205 2796 2209 2876
rect 2277 2796 2281 2876
rect 2285 2796 2289 2876
rect 2331 2836 2335 2876
rect 2417 2796 2421 2876
rect 2425 2796 2429 2876
rect 2471 2836 2475 2876
rect 2531 2836 2535 2876
rect 2553 2836 2557 2876
rect 2575 2796 2579 2876
rect 2636 2796 2640 2876
rect 2644 2796 2648 2876
rect 2666 2836 2670 2876
rect 2736 2796 2740 2876
rect 2744 2796 2748 2876
rect 2766 2836 2770 2876
rect 2831 2836 2835 2876
rect 2851 2836 2855 2876
rect 2915 2796 2919 2876
rect 2935 2836 2939 2876
rect 2949 2836 2953 2876
rect 2969 2836 2973 2876
rect 2981 2836 2985 2876
rect 3001 2836 3005 2876
rect 3047 2836 3051 2876
rect 3055 2836 3059 2876
rect 3075 2856 3079 2876
rect 3083 2856 3087 2876
rect 3105 2796 3109 2876
rect 3155 2796 3159 2876
rect 3175 2836 3179 2876
rect 3189 2836 3193 2876
rect 3209 2836 3213 2876
rect 3221 2836 3225 2876
rect 3241 2836 3245 2876
rect 3287 2836 3291 2876
rect 3295 2836 3299 2876
rect 3315 2856 3319 2876
rect 3323 2856 3327 2876
rect 3345 2796 3349 2876
rect 3405 2836 3409 2876
rect 3477 2796 3481 2876
rect 3485 2796 3489 2876
rect 3545 2796 3549 2876
rect 3595 2796 3599 2876
rect 3615 2836 3619 2876
rect 3629 2836 3633 2876
rect 3649 2836 3653 2876
rect 3661 2836 3665 2876
rect 3681 2836 3685 2876
rect 3727 2836 3731 2876
rect 3735 2836 3739 2876
rect 3755 2856 3759 2876
rect 3763 2856 3767 2876
rect 3785 2796 3789 2876
rect 3845 2796 3849 2876
rect 3865 2796 3869 2876
rect 3885 2796 3889 2876
rect 3905 2796 3909 2876
rect 3977 2796 3981 2876
rect 3985 2796 3989 2876
rect 4036 2796 4040 2876
rect 4044 2796 4048 2876
rect 4066 2836 4070 2876
rect 4150 2836 4154 2876
rect 4172 2796 4176 2876
rect 4180 2796 4184 2876
rect 4231 2796 4235 2876
rect 4239 2796 4243 2876
rect 4315 2796 4319 2876
rect 4335 2836 4339 2876
rect 4349 2836 4353 2876
rect 4369 2836 4373 2876
rect 4381 2836 4385 2876
rect 4401 2836 4405 2876
rect 4447 2836 4451 2876
rect 4455 2836 4459 2876
rect 4475 2856 4479 2876
rect 4483 2856 4487 2876
rect 4505 2796 4509 2876
rect 4556 2796 4560 2876
rect 4564 2796 4568 2876
rect 4586 2836 4590 2876
rect 4651 2836 4655 2876
rect 4671 2836 4675 2876
rect 31 2424 35 2464
rect 51 2424 55 2464
rect 71 2424 75 2464
rect 131 2424 135 2504
rect 151 2424 155 2504
rect 171 2424 175 2504
rect 245 2424 249 2464
rect 301 2424 305 2504
rect 323 2424 327 2464
rect 345 2424 349 2464
rect 405 2424 409 2504
rect 425 2424 429 2504
rect 445 2424 449 2504
rect 505 2424 509 2464
rect 525 2424 529 2464
rect 545 2424 549 2464
rect 610 2424 614 2464
rect 632 2424 636 2504
rect 640 2424 644 2504
rect 705 2424 709 2504
rect 765 2424 769 2464
rect 785 2424 789 2464
rect 845 2424 849 2464
rect 865 2424 869 2464
rect 885 2424 889 2464
rect 950 2424 954 2464
rect 972 2424 976 2504
rect 980 2424 984 2504
rect 1031 2424 1035 2464
rect 1051 2424 1055 2464
rect 1125 2424 1129 2464
rect 1145 2424 1149 2464
rect 1165 2424 1169 2464
rect 1225 2424 1229 2464
rect 1290 2424 1294 2464
rect 1312 2424 1316 2504
rect 1320 2424 1324 2504
rect 1371 2424 1375 2464
rect 1391 2424 1395 2464
rect 1451 2424 1455 2504
rect 1525 2424 1529 2464
rect 1545 2424 1549 2464
rect 1595 2424 1599 2504
rect 1615 2424 1619 2464
rect 1629 2424 1633 2464
rect 1649 2424 1653 2464
rect 1661 2424 1665 2464
rect 1681 2424 1685 2464
rect 1727 2424 1731 2464
rect 1735 2424 1739 2464
rect 1755 2424 1759 2444
rect 1763 2424 1767 2444
rect 1785 2424 1789 2504
rect 1831 2424 1835 2464
rect 1851 2424 1855 2464
rect 1911 2424 1915 2464
rect 1931 2424 1935 2464
rect 1991 2424 1995 2464
rect 2011 2424 2015 2464
rect 2031 2424 2035 2464
rect 2091 2424 2095 2504
rect 2099 2424 2103 2504
rect 2185 2424 2189 2464
rect 2257 2424 2261 2504
rect 2265 2424 2269 2504
rect 2325 2424 2329 2464
rect 2390 2424 2394 2464
rect 2412 2424 2416 2504
rect 2420 2424 2424 2504
rect 2471 2424 2475 2504
rect 2479 2424 2483 2504
rect 2551 2424 2555 2464
rect 2573 2424 2577 2464
rect 2595 2424 2599 2504
rect 2656 2424 2660 2504
rect 2664 2424 2668 2504
rect 2686 2424 2690 2464
rect 2765 2424 2769 2464
rect 2785 2424 2789 2464
rect 2831 2424 2835 2504
rect 2841 2424 2845 2504
rect 2861 2424 2865 2504
rect 2931 2424 2935 2464
rect 2951 2424 2955 2464
rect 3011 2424 3015 2464
rect 3033 2424 3037 2504
rect 3096 2424 3100 2504
rect 3104 2424 3108 2504
rect 3126 2424 3130 2464
rect 3203 2424 3207 2504
rect 3225 2424 3229 2464
rect 3285 2424 3289 2464
rect 3305 2424 3309 2464
rect 3351 2424 3355 2504
rect 3371 2424 3375 2504
rect 3391 2424 3395 2504
rect 3411 2424 3415 2504
rect 3471 2424 3475 2464
rect 3493 2424 3497 2504
rect 3563 2424 3567 2504
rect 3585 2424 3589 2464
rect 3635 2424 3639 2504
rect 3655 2424 3659 2464
rect 3669 2424 3673 2464
rect 3689 2424 3693 2464
rect 3701 2424 3705 2464
rect 3721 2424 3725 2464
rect 3767 2424 3771 2464
rect 3775 2424 3779 2464
rect 3795 2424 3799 2444
rect 3803 2424 3807 2444
rect 3825 2424 3829 2504
rect 3885 2424 3889 2504
rect 3905 2424 3909 2504
rect 3925 2424 3929 2504
rect 3971 2424 3975 2504
rect 3979 2424 3983 2504
rect 4051 2424 4055 2504
rect 4071 2424 4075 2504
rect 4091 2424 4095 2504
rect 4111 2424 4115 2504
rect 4131 2424 4135 2504
rect 4151 2424 4155 2504
rect 4171 2424 4175 2504
rect 4191 2424 4195 2504
rect 4255 2424 4259 2504
rect 4275 2424 4279 2464
rect 4289 2424 4293 2464
rect 4309 2424 4313 2464
rect 4321 2424 4325 2464
rect 4341 2424 4345 2464
rect 4387 2424 4391 2464
rect 4395 2424 4399 2464
rect 4415 2424 4419 2444
rect 4423 2424 4427 2444
rect 4445 2424 4449 2504
rect 4496 2424 4500 2504
rect 4504 2424 4508 2504
rect 4526 2424 4530 2464
rect 4591 2424 4595 2464
rect 4611 2424 4615 2464
rect 4671 2424 4675 2464
rect 4691 2424 4695 2464
rect 45 2356 49 2396
rect 65 2356 69 2396
rect 85 2356 89 2396
rect 150 2356 154 2396
rect 172 2316 176 2396
rect 180 2316 184 2396
rect 236 2316 240 2396
rect 244 2316 248 2396
rect 266 2356 270 2396
rect 331 2356 335 2396
rect 351 2356 355 2396
rect 371 2356 375 2396
rect 431 2316 435 2396
rect 451 2316 455 2396
rect 471 2316 475 2396
rect 536 2316 540 2396
rect 544 2316 548 2396
rect 566 2356 570 2396
rect 645 2316 649 2396
rect 665 2316 669 2396
rect 685 2316 689 2396
rect 731 2356 735 2396
rect 801 2316 805 2396
rect 823 2356 827 2396
rect 845 2356 849 2396
rect 891 2356 895 2396
rect 911 2356 915 2396
rect 971 2356 975 2396
rect 993 2356 997 2396
rect 1015 2316 1019 2396
rect 1090 2356 1094 2396
rect 1112 2316 1116 2396
rect 1120 2316 1124 2396
rect 1190 2356 1194 2396
rect 1212 2316 1216 2396
rect 1220 2316 1224 2396
rect 1275 2316 1279 2396
rect 1295 2356 1299 2396
rect 1309 2356 1313 2396
rect 1329 2356 1333 2396
rect 1341 2356 1345 2396
rect 1361 2356 1365 2396
rect 1407 2356 1411 2396
rect 1415 2356 1419 2396
rect 1435 2376 1439 2396
rect 1443 2376 1447 2396
rect 1465 2316 1469 2396
rect 1530 2356 1534 2396
rect 1552 2316 1556 2396
rect 1560 2316 1564 2396
rect 1615 2316 1619 2396
rect 1635 2356 1639 2396
rect 1649 2356 1653 2396
rect 1669 2356 1673 2396
rect 1681 2356 1685 2396
rect 1701 2356 1705 2396
rect 1747 2356 1751 2396
rect 1755 2356 1759 2396
rect 1775 2376 1779 2396
rect 1783 2376 1787 2396
rect 1805 2316 1809 2396
rect 1865 2356 1869 2396
rect 1925 2356 1929 2396
rect 1976 2316 1980 2396
rect 1984 2316 1988 2396
rect 2006 2356 2010 2396
rect 2075 2316 2079 2396
rect 2095 2356 2099 2396
rect 2109 2356 2113 2396
rect 2129 2356 2133 2396
rect 2141 2356 2145 2396
rect 2161 2356 2165 2396
rect 2207 2356 2211 2396
rect 2215 2356 2219 2396
rect 2235 2376 2239 2396
rect 2243 2376 2247 2396
rect 2265 2316 2269 2396
rect 2325 2316 2329 2396
rect 2345 2316 2349 2396
rect 2365 2316 2369 2396
rect 2425 2316 2429 2396
rect 2445 2316 2449 2396
rect 2465 2316 2469 2396
rect 2511 2356 2515 2396
rect 2531 2356 2535 2396
rect 2551 2356 2555 2396
rect 2611 2356 2615 2396
rect 2633 2356 2637 2396
rect 2655 2316 2659 2396
rect 2711 2316 2715 2396
rect 2733 2376 2737 2396
rect 2741 2376 2745 2396
rect 2761 2356 2765 2396
rect 2769 2356 2773 2396
rect 2815 2356 2819 2396
rect 2835 2356 2839 2396
rect 2847 2356 2851 2396
rect 2867 2356 2871 2396
rect 2881 2356 2885 2396
rect 2901 2316 2905 2396
rect 2970 2356 2974 2396
rect 2992 2316 2996 2396
rect 3000 2316 3004 2396
rect 3070 2356 3074 2396
rect 3092 2316 3096 2396
rect 3100 2316 3104 2396
rect 3156 2316 3160 2396
rect 3164 2316 3168 2396
rect 3186 2356 3190 2396
rect 3251 2316 3255 2396
rect 3273 2376 3277 2396
rect 3281 2376 3285 2396
rect 3301 2356 3305 2396
rect 3309 2356 3313 2396
rect 3355 2356 3359 2396
rect 3375 2356 3379 2396
rect 3387 2356 3391 2396
rect 3407 2356 3411 2396
rect 3421 2356 3425 2396
rect 3441 2316 3445 2396
rect 3510 2356 3514 2396
rect 3532 2316 3536 2396
rect 3540 2316 3544 2396
rect 3617 2316 3621 2396
rect 3625 2316 3629 2396
rect 3671 2316 3675 2396
rect 3681 2316 3685 2396
rect 3701 2316 3705 2396
rect 3785 2356 3789 2396
rect 3805 2356 3809 2396
rect 3865 2316 3869 2396
rect 3885 2316 3889 2396
rect 3905 2316 3909 2396
rect 3925 2316 3929 2396
rect 3985 2316 3989 2396
rect 4005 2316 4009 2396
rect 4025 2316 4029 2396
rect 4045 2316 4049 2396
rect 4095 2316 4099 2396
rect 4115 2356 4119 2396
rect 4129 2356 4133 2396
rect 4149 2356 4153 2396
rect 4161 2356 4165 2396
rect 4181 2356 4185 2396
rect 4227 2356 4231 2396
rect 4235 2356 4239 2396
rect 4255 2376 4259 2396
rect 4263 2376 4267 2396
rect 4285 2316 4289 2396
rect 4331 2316 4335 2396
rect 4353 2376 4357 2396
rect 4361 2376 4365 2396
rect 4381 2356 4385 2396
rect 4389 2356 4393 2396
rect 4435 2356 4439 2396
rect 4455 2356 4459 2396
rect 4467 2356 4471 2396
rect 4487 2356 4491 2396
rect 4501 2356 4505 2396
rect 4521 2316 4525 2396
rect 4576 2316 4580 2396
rect 4584 2316 4588 2396
rect 4606 2356 4610 2396
rect 4671 2356 4675 2396
rect 4691 2356 4695 2396
rect 43 1944 47 2024
rect 65 1944 69 1984
rect 130 1944 134 1984
rect 152 1944 156 2024
rect 160 1944 164 2024
rect 225 1944 229 1984
rect 245 1944 249 1984
rect 265 1944 269 1984
rect 311 1944 315 2024
rect 331 1944 335 2024
rect 351 1944 355 2024
rect 411 1944 415 2024
rect 431 1944 435 2024
rect 451 1944 455 2024
rect 511 1944 515 1984
rect 531 1944 535 1984
rect 551 1944 555 1984
rect 611 1944 615 1984
rect 631 1944 635 1984
rect 651 1944 655 1984
rect 711 1944 715 2024
rect 731 1944 735 2024
rect 751 1944 755 2024
rect 830 1944 834 1984
rect 852 1944 856 2024
rect 860 1944 864 2024
rect 911 1944 915 1984
rect 931 1944 935 1984
rect 951 1944 955 1984
rect 1011 1944 1015 1984
rect 1031 1944 1035 1984
rect 1051 1944 1055 1984
rect 1111 1944 1115 1984
rect 1131 1944 1135 1984
rect 1151 1944 1155 1984
rect 1211 1944 1215 2024
rect 1231 1944 1235 2024
rect 1251 1944 1255 2024
rect 1311 1944 1315 2024
rect 1319 1944 1323 2024
rect 1405 1944 1409 1984
rect 1425 1944 1429 1984
rect 1485 1944 1489 1984
rect 1505 1944 1509 1984
rect 1551 1944 1555 1984
rect 1571 1944 1575 1984
rect 1650 1944 1654 1984
rect 1672 1944 1676 2024
rect 1680 1944 1684 2024
rect 1731 1944 1735 2024
rect 1751 1944 1755 2024
rect 1771 1944 1775 2024
rect 1831 1944 1835 2024
rect 1839 1944 1843 2024
rect 1930 1944 1934 1984
rect 1952 1944 1956 2024
rect 1960 1944 1964 2024
rect 2016 1944 2020 2024
rect 2024 1944 2028 2024
rect 2046 1944 2050 1984
rect 2130 1944 2134 1984
rect 2152 1944 2156 2024
rect 2160 1944 2164 2024
rect 2225 1944 2229 2024
rect 2245 1944 2249 2024
rect 2265 1944 2269 2024
rect 2285 1944 2289 2024
rect 2305 1944 2309 2024
rect 2325 1944 2329 2024
rect 2345 1944 2349 2024
rect 2365 1944 2369 2024
rect 2411 1944 2415 1984
rect 2431 1944 2435 1984
rect 2501 1944 2505 2024
rect 2523 1944 2527 1984
rect 2545 1944 2549 1984
rect 2591 1944 2595 2024
rect 2601 1944 2605 2024
rect 2621 1944 2625 2024
rect 2705 1944 2709 1984
rect 2725 1944 2729 1984
rect 2771 1944 2775 1984
rect 2791 1944 2795 1984
rect 2855 1944 2859 2024
rect 2875 1944 2879 1984
rect 2889 1944 2893 1984
rect 2909 1944 2913 1984
rect 2921 1944 2925 1984
rect 2941 1944 2945 1984
rect 2987 1944 2991 1984
rect 2995 1944 2999 1984
rect 3015 1944 3019 1964
rect 3023 1944 3027 1964
rect 3045 1944 3049 2024
rect 3105 1944 3109 2024
rect 3125 1944 3129 2024
rect 3145 1944 3149 2024
rect 3191 1944 3195 2024
rect 3199 1944 3203 2024
rect 3285 1944 3289 2024
rect 3305 1944 3309 2024
rect 3325 1944 3329 2024
rect 3345 1944 3349 2024
rect 3395 1944 3399 2024
rect 3415 1944 3419 1984
rect 3429 1944 3433 1984
rect 3449 1944 3453 1984
rect 3461 1944 3465 1984
rect 3481 1944 3485 1984
rect 3527 1944 3531 1984
rect 3535 1944 3539 1984
rect 3555 1944 3559 1964
rect 3563 1944 3567 1964
rect 3585 1944 3589 2024
rect 3636 1944 3640 2024
rect 3644 1944 3648 2024
rect 3666 1944 3670 1984
rect 3735 1944 3739 2024
rect 3755 1944 3759 1984
rect 3769 1944 3773 1984
rect 3789 1944 3793 1984
rect 3801 1944 3805 1984
rect 3821 1944 3825 1984
rect 3867 1944 3871 1984
rect 3875 1944 3879 1984
rect 3895 1944 3899 1964
rect 3903 1944 3907 1964
rect 3925 1944 3929 2024
rect 3971 1944 3975 2024
rect 3993 1944 3997 1964
rect 4001 1944 4005 1964
rect 4021 1944 4025 1984
rect 4029 1944 4033 1984
rect 4075 1944 4079 1984
rect 4095 1944 4099 1984
rect 4107 1944 4111 1984
rect 4127 1944 4131 1984
rect 4141 1944 4145 1984
rect 4161 1944 4165 2024
rect 4225 1944 4229 2024
rect 4245 1944 4249 2024
rect 4265 1944 4269 2024
rect 4285 1944 4289 2024
rect 4331 1944 4335 1984
rect 4417 1944 4421 2024
rect 4425 1944 4429 2024
rect 4497 1944 4501 2024
rect 4505 1944 4509 2024
rect 4551 1944 4555 2024
rect 4573 1944 4577 1964
rect 4581 1944 4585 1964
rect 4601 1944 4605 1984
rect 4609 1944 4613 1984
rect 4655 1944 4659 1984
rect 4675 1944 4679 1984
rect 4687 1944 4691 1984
rect 4707 1944 4711 1984
rect 4721 1944 4725 1984
rect 4741 1944 4745 2024
rect 45 1836 49 1916
rect 65 1836 69 1916
rect 85 1836 89 1916
rect 105 1836 109 1916
rect 156 1836 160 1916
rect 164 1836 168 1916
rect 186 1876 190 1916
rect 251 1876 255 1916
rect 271 1876 275 1916
rect 345 1876 349 1916
rect 365 1876 369 1916
rect 385 1876 389 1916
rect 431 1836 435 1916
rect 451 1836 455 1916
rect 471 1836 475 1916
rect 491 1836 495 1916
rect 551 1876 555 1916
rect 573 1876 577 1916
rect 595 1836 599 1916
rect 665 1836 669 1916
rect 711 1876 715 1916
rect 733 1836 737 1916
rect 810 1876 814 1916
rect 832 1836 836 1916
rect 840 1836 844 1916
rect 896 1836 900 1916
rect 904 1836 908 1916
rect 926 1876 930 1916
rect 991 1876 995 1916
rect 1011 1876 1015 1916
rect 1031 1876 1035 1916
rect 1091 1876 1095 1916
rect 1151 1876 1155 1916
rect 1171 1876 1175 1916
rect 1191 1876 1195 1916
rect 1251 1876 1255 1916
rect 1271 1876 1275 1916
rect 1291 1876 1295 1916
rect 1365 1876 1369 1916
rect 1425 1836 1429 1916
rect 1445 1836 1449 1916
rect 1465 1836 1469 1916
rect 1485 1836 1489 1916
rect 1531 1876 1535 1916
rect 1551 1876 1555 1916
rect 1571 1876 1575 1916
rect 1631 1876 1635 1916
rect 1705 1836 1709 1916
rect 1765 1876 1769 1916
rect 1785 1876 1789 1916
rect 1805 1876 1809 1916
rect 1851 1876 1855 1916
rect 1873 1876 1877 1916
rect 1895 1836 1899 1916
rect 1955 1836 1959 1916
rect 1975 1876 1979 1916
rect 1989 1876 1993 1916
rect 2009 1876 2013 1916
rect 2021 1876 2025 1916
rect 2041 1876 2045 1916
rect 2087 1876 2091 1916
rect 2095 1876 2099 1916
rect 2115 1896 2119 1916
rect 2123 1896 2127 1916
rect 2145 1836 2149 1916
rect 2217 1836 2221 1916
rect 2225 1836 2229 1916
rect 2271 1876 2275 1916
rect 2336 1836 2340 1916
rect 2344 1836 2348 1916
rect 2366 1876 2370 1916
rect 2431 1836 2435 1916
rect 2439 1836 2443 1916
rect 2511 1836 2515 1916
rect 2519 1836 2523 1916
rect 2596 1836 2600 1916
rect 2604 1836 2608 1916
rect 2626 1876 2630 1916
rect 2705 1876 2709 1916
rect 2725 1876 2729 1916
rect 2797 1836 2801 1916
rect 2805 1836 2809 1916
rect 2856 1836 2860 1916
rect 2864 1836 2868 1916
rect 2886 1876 2890 1916
rect 2951 1876 2955 1916
rect 3037 1836 3041 1916
rect 3045 1836 3049 1916
rect 3091 1836 3095 1916
rect 3113 1896 3117 1916
rect 3121 1896 3125 1916
rect 3141 1876 3145 1916
rect 3149 1876 3153 1916
rect 3195 1876 3199 1916
rect 3215 1876 3219 1916
rect 3227 1876 3231 1916
rect 3247 1876 3251 1916
rect 3261 1876 3265 1916
rect 3281 1836 3285 1916
rect 3336 1836 3340 1916
rect 3344 1836 3348 1916
rect 3366 1876 3370 1916
rect 3431 1876 3435 1916
rect 3451 1876 3455 1916
rect 3511 1836 3515 1916
rect 3533 1896 3537 1916
rect 3541 1896 3545 1916
rect 3561 1876 3565 1916
rect 3569 1876 3573 1916
rect 3615 1876 3619 1916
rect 3635 1876 3639 1916
rect 3647 1876 3651 1916
rect 3667 1876 3671 1916
rect 3681 1876 3685 1916
rect 3701 1836 3705 1916
rect 3751 1876 3755 1916
rect 3773 1836 3777 1916
rect 3845 1876 3849 1916
rect 3865 1876 3869 1916
rect 3930 1876 3934 1916
rect 3952 1836 3956 1916
rect 3960 1836 3964 1916
rect 4030 1876 4034 1916
rect 4052 1836 4056 1916
rect 4060 1836 4064 1916
rect 4111 1836 4115 1916
rect 4121 1836 4125 1916
rect 4141 1836 4145 1916
rect 4225 1876 4229 1916
rect 4271 1836 4275 1916
rect 4291 1836 4295 1916
rect 4311 1836 4315 1916
rect 4397 1836 4401 1916
rect 4405 1836 4409 1916
rect 4451 1836 4455 1916
rect 4473 1896 4477 1916
rect 4481 1896 4485 1916
rect 4501 1876 4505 1916
rect 4509 1876 4513 1916
rect 4555 1876 4559 1916
rect 4575 1876 4579 1916
rect 4587 1876 4591 1916
rect 4607 1876 4611 1916
rect 4621 1876 4625 1916
rect 4641 1836 4645 1916
rect 4705 1876 4709 1916
rect 4725 1876 4729 1916
rect 45 1464 49 1504
rect 105 1464 109 1544
rect 125 1464 129 1544
rect 145 1464 149 1544
rect 191 1464 195 1504
rect 211 1464 215 1504
rect 231 1464 235 1504
rect 291 1464 295 1504
rect 311 1464 315 1504
rect 390 1464 394 1504
rect 412 1464 416 1544
rect 420 1464 424 1544
rect 483 1464 487 1544
rect 505 1464 509 1504
rect 565 1464 569 1504
rect 611 1464 615 1504
rect 631 1464 635 1504
rect 651 1464 655 1504
rect 711 1464 715 1544
rect 731 1464 735 1544
rect 751 1464 755 1544
rect 811 1464 815 1504
rect 831 1464 835 1504
rect 851 1464 855 1504
rect 911 1464 915 1544
rect 931 1464 935 1544
rect 951 1464 955 1544
rect 1011 1464 1015 1504
rect 1031 1464 1035 1504
rect 1051 1464 1055 1504
rect 1130 1464 1134 1504
rect 1152 1464 1156 1544
rect 1160 1464 1164 1544
rect 1211 1464 1215 1504
rect 1231 1464 1235 1504
rect 1251 1464 1255 1504
rect 1311 1464 1315 1544
rect 1331 1464 1335 1544
rect 1351 1464 1355 1544
rect 1425 1464 1429 1504
rect 1471 1464 1475 1504
rect 1491 1464 1495 1504
rect 1511 1464 1515 1504
rect 1571 1464 1575 1544
rect 1591 1464 1595 1544
rect 1611 1464 1615 1544
rect 1671 1464 1675 1504
rect 1691 1464 1695 1504
rect 1711 1464 1715 1504
rect 1776 1464 1780 1544
rect 1784 1464 1788 1544
rect 1806 1464 1810 1504
rect 1885 1464 1889 1544
rect 1905 1464 1909 1544
rect 1925 1464 1929 1544
rect 1971 1464 1975 1504
rect 2031 1464 2035 1504
rect 2051 1464 2055 1504
rect 2071 1464 2075 1504
rect 2150 1464 2154 1504
rect 2172 1464 2176 1544
rect 2180 1464 2184 1544
rect 2231 1464 2235 1504
rect 2291 1464 2295 1544
rect 2313 1464 2317 1484
rect 2321 1464 2325 1484
rect 2341 1464 2345 1504
rect 2349 1464 2353 1504
rect 2395 1464 2399 1504
rect 2415 1464 2419 1504
rect 2427 1464 2431 1504
rect 2447 1464 2451 1504
rect 2461 1464 2465 1504
rect 2481 1464 2485 1544
rect 2550 1464 2554 1504
rect 2572 1464 2576 1544
rect 2580 1464 2584 1544
rect 2641 1464 2645 1544
rect 2663 1464 2667 1504
rect 2685 1464 2689 1504
rect 2731 1464 2735 1544
rect 2739 1464 2743 1544
rect 2811 1464 2815 1544
rect 2831 1464 2835 1544
rect 2851 1464 2855 1544
rect 2937 1464 2941 1544
rect 2945 1464 2949 1544
rect 3005 1464 3009 1504
rect 3065 1464 3069 1504
rect 3116 1464 3120 1544
rect 3124 1464 3128 1544
rect 3146 1464 3150 1504
rect 3211 1464 3215 1504
rect 3231 1464 3235 1504
rect 3305 1464 3309 1504
rect 3325 1464 3329 1504
rect 3390 1464 3394 1504
rect 3412 1464 3416 1544
rect 3420 1464 3424 1544
rect 3475 1464 3479 1544
rect 3495 1464 3499 1504
rect 3509 1464 3513 1504
rect 3529 1464 3533 1504
rect 3541 1464 3545 1504
rect 3561 1464 3565 1504
rect 3607 1464 3611 1504
rect 3615 1464 3619 1504
rect 3635 1464 3639 1484
rect 3643 1464 3647 1484
rect 3665 1464 3669 1544
rect 3711 1464 3715 1504
rect 3785 1464 3789 1504
rect 3850 1464 3854 1504
rect 3872 1464 3876 1544
rect 3880 1464 3884 1544
rect 3931 1464 3935 1544
rect 3939 1464 3943 1544
rect 4011 1464 4015 1544
rect 4019 1464 4023 1544
rect 4091 1464 4095 1504
rect 4151 1464 4155 1544
rect 4171 1464 4175 1544
rect 4191 1464 4195 1544
rect 4251 1464 4255 1544
rect 4259 1464 4263 1544
rect 4331 1464 4335 1544
rect 4351 1464 4355 1544
rect 4371 1464 4375 1544
rect 4431 1464 4435 1504
rect 4491 1464 4495 1504
rect 4565 1464 4569 1504
rect 4616 1464 4620 1544
rect 4624 1464 4628 1544
rect 4646 1464 4650 1504
rect 4711 1464 4715 1504
rect 4731 1464 4735 1504
rect 45 1356 49 1436
rect 65 1356 69 1436
rect 85 1356 89 1436
rect 131 1396 135 1436
rect 151 1396 155 1436
rect 171 1396 175 1436
rect 231 1396 235 1436
rect 251 1396 255 1436
rect 271 1396 275 1436
rect 345 1396 349 1436
rect 365 1396 369 1436
rect 416 1356 420 1436
rect 424 1356 428 1436
rect 446 1396 450 1436
rect 511 1356 515 1436
rect 531 1356 535 1436
rect 551 1356 555 1436
rect 616 1356 620 1436
rect 624 1356 628 1436
rect 646 1396 650 1436
rect 716 1356 720 1436
rect 724 1356 728 1436
rect 746 1396 750 1436
rect 811 1396 815 1436
rect 833 1396 837 1436
rect 855 1356 859 1436
rect 925 1396 929 1436
rect 945 1396 949 1436
rect 991 1396 995 1436
rect 1011 1396 1015 1436
rect 1085 1396 1089 1436
rect 1105 1396 1109 1436
rect 1125 1396 1129 1436
rect 1185 1396 1189 1436
rect 1241 1356 1245 1436
rect 1263 1396 1267 1436
rect 1285 1396 1289 1436
rect 1336 1356 1340 1436
rect 1344 1356 1348 1436
rect 1366 1396 1370 1436
rect 1450 1396 1454 1436
rect 1472 1356 1476 1436
rect 1480 1356 1484 1436
rect 1531 1396 1535 1436
rect 1551 1396 1555 1436
rect 1616 1356 1620 1436
rect 1624 1356 1628 1436
rect 1646 1396 1650 1436
rect 1711 1396 1715 1436
rect 1731 1396 1735 1436
rect 1791 1356 1795 1436
rect 1811 1356 1815 1436
rect 1831 1356 1835 1436
rect 1891 1396 1895 1436
rect 1911 1396 1915 1436
rect 1931 1396 1935 1436
rect 1996 1356 2000 1436
rect 2004 1356 2008 1436
rect 2026 1396 2030 1436
rect 2091 1396 2095 1436
rect 2151 1396 2155 1436
rect 2171 1396 2175 1436
rect 2191 1396 2195 1436
rect 2251 1396 2255 1436
rect 2271 1396 2275 1436
rect 2331 1356 2335 1436
rect 2341 1356 2345 1436
rect 2361 1356 2365 1436
rect 2445 1396 2449 1436
rect 2465 1396 2469 1436
rect 2511 1396 2515 1436
rect 2583 1356 2587 1436
rect 2605 1396 2609 1436
rect 2656 1356 2660 1436
rect 2664 1356 2668 1436
rect 2686 1396 2690 1436
rect 2775 1356 2779 1436
rect 2785 1356 2789 1436
rect 2815 1356 2819 1436
rect 2825 1356 2829 1436
rect 2875 1356 2879 1436
rect 2895 1396 2899 1436
rect 2909 1396 2913 1436
rect 2929 1396 2933 1436
rect 2941 1396 2945 1436
rect 2961 1396 2965 1436
rect 3007 1396 3011 1436
rect 3015 1396 3019 1436
rect 3035 1416 3039 1436
rect 3043 1416 3047 1436
rect 3065 1356 3069 1436
rect 3137 1356 3141 1436
rect 3145 1356 3149 1436
rect 3205 1356 3209 1436
rect 3225 1356 3229 1436
rect 3245 1356 3249 1436
rect 3295 1356 3299 1436
rect 3315 1396 3319 1436
rect 3329 1396 3333 1436
rect 3349 1396 3353 1436
rect 3361 1396 3365 1436
rect 3381 1396 3385 1436
rect 3427 1396 3431 1436
rect 3435 1396 3439 1436
rect 3455 1416 3459 1436
rect 3463 1416 3467 1436
rect 3485 1356 3489 1436
rect 3545 1396 3549 1436
rect 3617 1356 3621 1436
rect 3625 1356 3629 1436
rect 3697 1356 3701 1436
rect 3705 1356 3709 1436
rect 3751 1396 3755 1436
rect 3811 1356 3815 1436
rect 3833 1416 3837 1436
rect 3841 1416 3845 1436
rect 3861 1396 3865 1436
rect 3869 1396 3873 1436
rect 3915 1396 3919 1436
rect 3935 1396 3939 1436
rect 3947 1396 3951 1436
rect 3967 1396 3971 1436
rect 3981 1396 3985 1436
rect 4001 1356 4005 1436
rect 4056 1356 4060 1436
rect 4064 1356 4068 1436
rect 4086 1396 4090 1436
rect 4151 1396 4155 1436
rect 4171 1396 4175 1436
rect 4243 1356 4247 1436
rect 4265 1396 4269 1436
rect 4325 1396 4329 1436
rect 4345 1396 4349 1436
rect 4410 1396 4414 1436
rect 4432 1356 4436 1436
rect 4440 1356 4444 1436
rect 4510 1396 4514 1436
rect 4532 1356 4536 1436
rect 4540 1356 4544 1436
rect 4591 1356 4595 1436
rect 4599 1356 4603 1436
rect 4671 1396 4675 1436
rect 4745 1396 4749 1436
rect 50 984 54 1024
rect 72 984 76 1064
rect 80 984 84 1064
rect 136 984 140 1064
rect 144 984 148 1064
rect 166 984 170 1024
rect 231 984 235 1024
rect 251 984 255 1024
rect 271 984 275 1024
rect 331 984 335 1064
rect 351 984 355 1064
rect 371 984 375 1064
rect 431 984 435 1024
rect 451 984 455 1024
rect 471 984 475 1024
rect 531 984 535 1064
rect 551 984 555 1064
rect 571 984 575 1064
rect 645 984 649 1024
rect 665 984 669 1024
rect 721 984 725 1064
rect 743 984 747 1024
rect 765 984 769 1024
rect 825 984 829 1024
rect 845 984 849 1024
rect 865 984 869 1024
rect 930 984 934 1024
rect 952 984 956 1064
rect 960 984 964 1064
rect 1016 984 1020 1064
rect 1024 984 1028 1064
rect 1046 984 1050 1024
rect 1130 984 1134 1024
rect 1152 984 1156 1064
rect 1160 984 1164 1064
rect 1225 984 1229 1024
rect 1245 984 1249 1024
rect 1301 984 1305 1064
rect 1323 984 1327 1024
rect 1345 984 1349 1024
rect 1391 984 1395 1024
rect 1411 984 1415 1024
rect 1485 984 1489 1064
rect 1545 984 1549 1024
rect 1565 984 1569 1024
rect 1625 984 1629 1024
rect 1645 984 1649 1024
rect 1691 984 1695 1024
rect 1711 984 1715 1024
rect 1731 984 1735 1024
rect 1805 984 1809 1024
rect 1825 984 1829 1024
rect 1871 984 1875 1024
rect 1891 984 1895 1024
rect 1911 984 1915 1024
rect 1971 984 1975 1024
rect 1991 984 1995 1024
rect 2065 984 2069 1064
rect 2085 984 2089 1064
rect 2105 984 2109 1064
rect 2125 984 2129 1064
rect 2185 984 2189 1024
rect 2205 984 2209 1024
rect 2225 984 2229 1024
rect 2285 984 2289 1024
rect 2305 984 2309 1024
rect 2351 984 2355 1064
rect 2371 984 2375 1064
rect 2391 984 2395 1064
rect 2465 984 2469 1024
rect 2525 984 2529 1024
rect 2545 984 2549 1024
rect 2615 984 2619 1064
rect 2625 984 2629 1064
rect 2655 984 2659 1064
rect 2665 984 2669 1064
rect 2711 984 2715 1024
rect 2733 984 2737 1064
rect 2795 984 2799 1064
rect 2815 984 2819 1024
rect 2829 984 2833 1024
rect 2849 984 2853 1024
rect 2861 984 2865 1024
rect 2881 984 2885 1024
rect 2927 984 2931 1024
rect 2935 984 2939 1024
rect 2955 984 2959 1004
rect 2963 984 2967 1004
rect 2985 984 2989 1064
rect 3031 984 3035 1024
rect 3051 984 3055 1024
rect 3130 984 3134 1024
rect 3152 984 3156 1064
rect 3160 984 3164 1064
rect 3211 984 3215 1064
rect 3231 984 3235 1064
rect 3251 984 3255 1064
rect 3271 984 3275 1064
rect 3343 984 3347 1064
rect 3365 984 3369 1024
rect 3411 984 3415 1024
rect 3433 984 3437 1064
rect 3491 984 3495 1064
rect 3511 984 3515 1064
rect 3531 984 3535 1064
rect 3551 984 3555 1064
rect 3571 984 3575 1064
rect 3591 984 3595 1064
rect 3611 984 3615 1064
rect 3631 984 3635 1064
rect 3691 984 3695 1064
rect 3711 984 3715 1064
rect 3731 984 3735 1064
rect 3751 984 3755 1064
rect 3771 984 3775 1064
rect 3791 984 3795 1064
rect 3811 984 3815 1064
rect 3831 984 3835 1064
rect 3891 984 3895 1024
rect 3913 984 3917 1064
rect 3971 984 3975 1024
rect 3991 984 3995 1024
rect 4051 984 4055 1064
rect 4073 984 4077 1004
rect 4081 984 4085 1004
rect 4101 984 4105 1024
rect 4109 984 4113 1024
rect 4155 984 4159 1024
rect 4175 984 4179 1024
rect 4187 984 4191 1024
rect 4207 984 4211 1024
rect 4221 984 4225 1024
rect 4241 984 4245 1064
rect 4291 984 4295 1024
rect 4311 984 4315 1024
rect 4376 984 4380 1064
rect 4384 984 4388 1064
rect 4406 984 4410 1024
rect 4485 984 4489 1024
rect 4505 984 4509 1024
rect 4556 984 4560 1064
rect 4564 984 4568 1064
rect 4586 984 4590 1024
rect 4651 984 4655 1024
rect 4671 984 4675 1024
rect 4691 984 4695 1024
rect 45 916 49 956
rect 65 916 69 956
rect 121 876 125 956
rect 143 916 147 956
rect 165 916 169 956
rect 230 916 234 956
rect 252 876 256 956
rect 260 876 264 956
rect 325 876 329 956
rect 345 876 349 956
rect 365 876 369 956
rect 385 876 389 956
rect 443 876 447 956
rect 465 916 469 956
rect 511 916 515 956
rect 585 916 589 956
rect 645 876 649 956
rect 665 876 669 956
rect 685 876 689 956
rect 731 916 735 956
rect 751 916 755 956
rect 771 916 775 956
rect 841 876 845 956
rect 863 916 867 956
rect 885 916 889 956
rect 931 916 935 956
rect 951 916 955 956
rect 1025 916 1029 956
rect 1045 916 1049 956
rect 1065 916 1069 956
rect 1116 876 1120 956
rect 1124 876 1128 956
rect 1146 916 1150 956
rect 1225 916 1229 956
rect 1245 916 1249 956
rect 1265 916 1269 956
rect 1311 916 1315 956
rect 1376 876 1380 956
rect 1384 876 1388 956
rect 1406 916 1410 956
rect 1485 916 1489 956
rect 1505 916 1509 956
rect 1551 916 1555 956
rect 1571 916 1575 956
rect 1650 916 1654 956
rect 1672 876 1676 956
rect 1680 876 1684 956
rect 1731 916 1735 956
rect 1753 916 1757 956
rect 1775 876 1779 956
rect 1845 916 1849 956
rect 1905 916 1909 956
rect 1925 916 1929 956
rect 1971 916 1975 956
rect 2045 916 2049 956
rect 2065 916 2069 956
rect 2085 916 2089 956
rect 2131 916 2135 956
rect 2196 876 2200 956
rect 2204 876 2208 956
rect 2226 916 2230 956
rect 2305 876 2309 956
rect 2325 876 2329 956
rect 2345 876 2349 956
rect 2391 916 2395 956
rect 2451 916 2455 956
rect 2471 916 2475 956
rect 2491 916 2495 956
rect 2565 916 2569 956
rect 2585 916 2589 956
rect 2605 916 2609 956
rect 2651 876 2655 956
rect 2671 876 2675 956
rect 2691 876 2695 956
rect 2765 916 2769 956
rect 2785 916 2789 956
rect 2855 876 2859 956
rect 2865 876 2869 956
rect 2895 876 2899 956
rect 2905 876 2909 956
rect 2965 916 2969 956
rect 3037 876 3041 956
rect 3045 876 3049 956
rect 3117 876 3121 956
rect 3125 876 3129 956
rect 3171 916 3175 956
rect 3236 876 3240 956
rect 3244 876 3248 956
rect 3266 916 3270 956
rect 3331 916 3335 956
rect 3351 916 3355 956
rect 3411 876 3415 956
rect 3433 936 3437 956
rect 3441 936 3445 956
rect 3461 916 3465 956
rect 3469 916 3473 956
rect 3515 916 3519 956
rect 3535 916 3539 956
rect 3547 916 3551 956
rect 3567 916 3571 956
rect 3581 916 3585 956
rect 3601 876 3605 956
rect 3651 916 3655 956
rect 3673 876 3677 956
rect 3735 876 3739 956
rect 3755 916 3759 956
rect 3769 916 3773 956
rect 3789 916 3793 956
rect 3801 916 3805 956
rect 3821 916 3825 956
rect 3867 916 3871 956
rect 3875 916 3879 956
rect 3895 936 3899 956
rect 3903 936 3907 956
rect 3925 876 3929 956
rect 3990 916 3994 956
rect 4012 876 4016 956
rect 4020 876 4024 956
rect 4071 876 4075 956
rect 4093 936 4097 956
rect 4101 936 4105 956
rect 4121 916 4125 956
rect 4129 916 4133 956
rect 4175 916 4179 956
rect 4195 916 4199 956
rect 4207 916 4211 956
rect 4227 916 4231 956
rect 4241 916 4245 956
rect 4261 876 4265 956
rect 4315 876 4319 956
rect 4335 916 4339 956
rect 4349 916 4353 956
rect 4369 916 4373 956
rect 4381 916 4385 956
rect 4401 916 4405 956
rect 4447 916 4451 956
rect 4455 916 4459 956
rect 4475 936 4479 956
rect 4483 936 4487 956
rect 4505 876 4509 956
rect 4556 876 4560 956
rect 4564 876 4568 956
rect 4586 916 4590 956
rect 4656 876 4660 956
rect 4664 876 4668 956
rect 4686 916 4690 956
rect 57 504 61 584
rect 65 504 69 584
rect 125 504 129 584
rect 145 504 149 584
rect 165 504 169 584
rect 211 504 215 544
rect 285 504 289 584
rect 305 504 309 584
rect 325 504 329 584
rect 371 504 375 544
rect 391 504 395 544
rect 411 504 415 544
rect 490 504 494 544
rect 512 504 516 584
rect 520 504 524 584
rect 583 504 587 584
rect 605 504 609 544
rect 670 504 674 544
rect 692 504 696 584
rect 700 504 704 584
rect 763 504 767 584
rect 785 504 789 544
rect 831 504 835 544
rect 853 504 857 544
rect 875 504 879 584
rect 936 504 940 584
rect 944 504 948 584
rect 966 504 970 544
rect 1050 504 1054 544
rect 1072 504 1076 584
rect 1080 504 1084 584
rect 1145 504 1149 584
rect 1191 504 1195 584
rect 1211 504 1215 584
rect 1231 504 1235 584
rect 1305 504 1309 544
rect 1356 504 1360 584
rect 1364 504 1368 584
rect 1386 504 1390 544
rect 1456 504 1460 584
rect 1464 504 1468 584
rect 1486 504 1490 544
rect 1565 504 1569 584
rect 1585 504 1589 584
rect 1605 504 1609 584
rect 1651 504 1655 584
rect 1671 504 1675 584
rect 1691 504 1695 584
rect 1751 504 1755 544
rect 1771 504 1775 544
rect 1791 504 1795 544
rect 1856 504 1860 584
rect 1864 504 1868 584
rect 1886 504 1890 544
rect 1965 504 1969 584
rect 1985 504 1989 584
rect 2005 504 2009 584
rect 2056 504 2060 584
rect 2064 504 2068 584
rect 2086 504 2090 544
rect 2165 504 2169 544
rect 2185 504 2189 544
rect 2205 504 2209 544
rect 2270 504 2274 544
rect 2292 504 2296 584
rect 2300 504 2304 584
rect 2356 504 2360 584
rect 2364 504 2368 584
rect 2386 504 2390 544
rect 2451 504 2455 544
rect 2471 504 2475 544
rect 2491 504 2495 544
rect 2551 504 2555 544
rect 2571 504 2575 544
rect 2591 504 2595 544
rect 2665 504 2669 544
rect 2711 504 2715 544
rect 2731 504 2735 544
rect 2751 504 2755 544
rect 2815 504 2819 584
rect 2835 504 2839 544
rect 2849 504 2853 544
rect 2869 504 2873 544
rect 2881 504 2885 544
rect 2901 504 2905 544
rect 2947 504 2951 544
rect 2955 504 2959 544
rect 2975 504 2979 524
rect 2983 504 2987 524
rect 3005 504 3009 584
rect 3056 504 3060 584
rect 3064 504 3068 584
rect 3086 504 3090 544
rect 3151 504 3155 544
rect 3211 504 3215 544
rect 3271 504 3275 544
rect 3291 504 3295 544
rect 3311 504 3315 544
rect 3385 504 3389 544
rect 3445 504 3449 544
rect 3465 504 3469 544
rect 3530 504 3534 544
rect 3552 504 3556 584
rect 3560 504 3564 584
rect 3615 504 3619 584
rect 3635 504 3639 544
rect 3649 504 3653 544
rect 3669 504 3673 544
rect 3681 504 3685 544
rect 3701 504 3705 544
rect 3747 504 3751 544
rect 3755 504 3759 544
rect 3775 504 3779 524
rect 3783 504 3787 524
rect 3805 504 3809 584
rect 3856 504 3860 584
rect 3864 504 3868 584
rect 3886 504 3890 544
rect 3965 504 3969 544
rect 3985 504 3989 544
rect 4031 504 4035 584
rect 4053 504 4057 524
rect 4061 504 4065 524
rect 4081 504 4085 544
rect 4089 504 4093 544
rect 4135 504 4139 544
rect 4155 504 4159 544
rect 4167 504 4171 544
rect 4187 504 4191 544
rect 4201 504 4205 544
rect 4221 504 4225 584
rect 4271 504 4275 544
rect 4291 504 4295 544
rect 4351 504 4355 544
rect 4371 504 4375 544
rect 4450 504 4454 544
rect 4472 504 4476 584
rect 4480 504 4484 584
rect 4535 504 4539 584
rect 4555 504 4559 544
rect 4569 504 4573 544
rect 4589 504 4593 544
rect 4601 504 4605 544
rect 4621 504 4625 544
rect 4667 504 4671 544
rect 4675 504 4679 544
rect 4695 504 4699 524
rect 4703 504 4707 524
rect 4725 504 4729 584
rect 31 436 35 476
rect 51 436 55 476
rect 111 436 115 476
rect 131 436 135 476
rect 205 436 209 476
rect 225 436 229 476
rect 285 436 289 476
rect 305 436 309 476
rect 361 396 365 476
rect 383 436 387 476
rect 405 436 409 476
rect 465 436 469 476
rect 485 436 489 476
rect 545 436 549 476
rect 565 436 569 476
rect 585 436 589 476
rect 645 396 649 476
rect 665 396 669 476
rect 685 396 689 476
rect 705 396 709 476
rect 777 396 781 476
rect 785 396 789 476
rect 845 436 849 476
rect 865 436 869 476
rect 911 436 915 476
rect 931 436 935 476
rect 1005 436 1009 476
rect 1025 436 1029 476
rect 1085 436 1089 476
rect 1105 436 1109 476
rect 1165 396 1169 476
rect 1185 396 1189 476
rect 1205 396 1209 476
rect 1225 396 1229 476
rect 1276 396 1280 476
rect 1284 396 1288 476
rect 1306 436 1310 476
rect 1397 396 1401 476
rect 1405 396 1409 476
rect 1456 396 1460 476
rect 1464 396 1468 476
rect 1486 436 1490 476
rect 1551 436 1555 476
rect 1625 396 1629 476
rect 1645 396 1649 476
rect 1665 396 1669 476
rect 1711 436 1715 476
rect 1771 436 1775 476
rect 1791 436 1795 476
rect 1811 436 1815 476
rect 1871 396 1875 476
rect 1891 396 1895 476
rect 1911 396 1915 476
rect 1971 436 1975 476
rect 1991 436 1995 476
rect 2051 436 2055 476
rect 2071 436 2075 476
rect 2131 436 2135 476
rect 2151 436 2155 476
rect 2237 396 2241 476
rect 2245 396 2249 476
rect 2305 436 2309 476
rect 2325 436 2329 476
rect 2371 396 2375 476
rect 2379 396 2383 476
rect 2451 436 2455 476
rect 2471 436 2475 476
rect 2491 436 2495 476
rect 2565 436 2569 476
rect 2625 436 2629 476
rect 2645 436 2649 476
rect 2665 436 2669 476
rect 2711 396 2715 476
rect 2731 396 2735 476
rect 2751 396 2755 476
rect 2811 396 2815 476
rect 2819 396 2823 476
rect 2905 436 2909 476
rect 2925 436 2929 476
rect 2990 436 2994 476
rect 3012 396 3016 476
rect 3020 396 3024 476
rect 3090 436 3094 476
rect 3112 396 3116 476
rect 3120 396 3124 476
rect 3197 396 3201 476
rect 3205 396 3209 476
rect 3265 436 3269 476
rect 3330 436 3334 476
rect 3352 396 3356 476
rect 3360 396 3364 476
rect 3425 396 3429 476
rect 3445 396 3449 476
rect 3465 396 3469 476
rect 3537 396 3541 476
rect 3545 396 3549 476
rect 3591 396 3595 476
rect 3601 396 3605 476
rect 3621 396 3625 476
rect 3691 436 3695 476
rect 3711 436 3715 476
rect 3771 436 3775 476
rect 3791 436 3795 476
rect 3870 436 3874 476
rect 3892 396 3896 476
rect 3900 396 3904 476
rect 3965 436 3969 476
rect 4025 436 4029 476
rect 4071 396 4075 476
rect 4093 456 4097 476
rect 4101 456 4105 476
rect 4121 436 4125 476
rect 4129 436 4133 476
rect 4175 436 4179 476
rect 4195 436 4199 476
rect 4207 436 4211 476
rect 4227 436 4231 476
rect 4241 436 4245 476
rect 4261 396 4265 476
rect 4325 436 4329 476
rect 4345 436 4349 476
rect 4410 436 4414 476
rect 4432 396 4436 476
rect 4440 396 4444 476
rect 4505 436 4509 476
rect 4551 396 4555 476
rect 4573 456 4577 476
rect 4581 456 4585 476
rect 4601 436 4605 476
rect 4609 436 4613 476
rect 4655 436 4659 476
rect 4675 436 4679 476
rect 4687 436 4691 476
rect 4707 436 4711 476
rect 4721 436 4725 476
rect 4741 396 4745 476
rect 45 24 49 64
rect 65 24 69 64
rect 85 24 89 64
rect 131 24 135 104
rect 151 24 155 104
rect 171 24 175 104
rect 250 24 254 64
rect 272 24 276 104
rect 280 24 284 104
rect 336 24 340 104
rect 344 24 348 104
rect 366 24 370 64
rect 445 24 449 64
rect 465 24 469 64
rect 485 24 489 64
rect 531 24 535 64
rect 551 24 555 64
rect 571 24 575 64
rect 631 24 635 104
rect 651 24 655 104
rect 671 24 675 104
rect 745 24 749 104
rect 765 24 769 104
rect 785 24 789 104
rect 831 24 835 64
rect 910 24 914 64
rect 932 24 936 104
rect 940 24 944 104
rect 1005 24 1009 64
rect 1056 24 1060 104
rect 1064 24 1068 104
rect 1086 24 1090 64
rect 1156 24 1160 104
rect 1164 24 1168 104
rect 1186 24 1190 64
rect 1251 24 1255 64
rect 1271 24 1275 64
rect 1291 24 1295 64
rect 1351 24 1355 64
rect 1371 24 1375 64
rect 1391 24 1395 64
rect 1465 24 1469 104
rect 1485 24 1489 104
rect 1505 24 1509 104
rect 1551 24 1555 64
rect 1571 24 1575 64
rect 1591 24 1595 64
rect 1665 24 1669 104
rect 1685 24 1689 104
rect 1705 24 1709 104
rect 1751 24 1755 64
rect 1771 24 1775 64
rect 1791 24 1795 64
rect 1851 24 1855 64
rect 1871 24 1875 64
rect 1931 24 1935 64
rect 1953 24 1957 104
rect 2021 24 2025 104
rect 2043 24 2047 64
rect 2065 24 2069 64
rect 2111 24 2115 64
rect 2133 24 2137 104
rect 2191 24 2195 64
rect 2211 24 2215 64
rect 2231 24 2235 64
rect 2291 24 2295 104
rect 2311 24 2315 104
rect 2331 24 2335 104
rect 2351 24 2355 104
rect 2416 24 2420 104
rect 2424 24 2428 104
rect 2446 24 2450 64
rect 2525 24 2529 104
rect 2545 24 2549 104
rect 2565 24 2569 104
rect 2616 24 2620 104
rect 2624 24 2628 104
rect 2646 24 2650 64
rect 2711 24 2715 64
rect 2771 24 2775 64
rect 2791 24 2795 64
rect 2811 24 2815 64
rect 2871 24 2875 64
rect 2935 24 2939 104
rect 2955 24 2959 64
rect 2969 24 2973 64
rect 2989 24 2993 64
rect 3001 24 3005 64
rect 3021 24 3025 64
rect 3067 24 3071 64
rect 3075 24 3079 64
rect 3095 24 3099 44
rect 3103 24 3107 44
rect 3125 24 3129 104
rect 3171 24 3175 64
rect 3245 24 3249 64
rect 3295 24 3299 104
rect 3315 24 3319 64
rect 3329 24 3333 64
rect 3349 24 3353 64
rect 3361 24 3365 64
rect 3381 24 3385 64
rect 3427 24 3431 64
rect 3435 24 3439 64
rect 3455 24 3459 44
rect 3463 24 3467 44
rect 3485 24 3489 104
rect 3557 24 3561 104
rect 3565 24 3569 104
rect 3611 24 3615 104
rect 3633 24 3637 44
rect 3641 24 3645 44
rect 3661 24 3665 64
rect 3669 24 3673 64
rect 3715 24 3719 64
rect 3735 24 3739 64
rect 3747 24 3751 64
rect 3767 24 3771 64
rect 3781 24 3785 64
rect 3801 24 3805 104
rect 3851 24 3855 64
rect 3916 24 3920 104
rect 3924 24 3928 104
rect 3946 24 3950 64
rect 4011 24 4015 104
rect 4019 24 4023 104
rect 4091 24 4095 104
rect 4099 24 4103 104
rect 4197 24 4201 104
rect 4205 24 4209 104
rect 4256 24 4260 104
rect 4264 24 4268 104
rect 4286 24 4290 64
rect 4365 24 4369 64
rect 4385 24 4389 64
rect 4445 24 4449 64
rect 4491 24 4495 104
rect 4499 24 4503 104
rect 4571 24 4575 64
rect 4591 24 4595 64
rect 4665 24 4669 64
rect 4711 24 4715 64
rect 4731 24 4735 64
<< ndiffusion >>
rect 50 4536 52 4556
rect 56 4536 60 4556
rect 72 4516 74 4556
rect 78 4516 82 4556
rect 86 4516 88 4556
rect 166 4498 168 4556
rect 154 4496 168 4498
rect 172 4496 176 4556
rect 180 4496 184 4556
rect 188 4496 190 4556
rect 230 4496 232 4556
rect 236 4496 240 4556
rect 244 4496 248 4556
rect 252 4498 254 4556
rect 252 4496 266 4498
rect 366 4498 368 4556
rect 354 4496 368 4498
rect 372 4496 376 4556
rect 380 4496 384 4556
rect 388 4496 390 4556
rect 432 4516 434 4556
rect 438 4516 442 4556
rect 446 4516 448 4556
rect 460 4536 464 4556
rect 468 4536 470 4556
rect 529 4516 531 4556
rect 535 4528 537 4556
rect 549 4528 551 4556
rect 535 4516 551 4528
rect 555 4516 557 4556
rect 569 4516 571 4556
rect 575 4516 577 4556
rect 629 4516 631 4556
rect 635 4528 637 4556
rect 649 4528 651 4556
rect 635 4516 651 4528
rect 655 4516 657 4556
rect 669 4516 671 4556
rect 675 4516 677 4556
rect 766 4498 768 4556
rect 754 4496 768 4498
rect 772 4496 776 4556
rect 780 4496 784 4556
rect 788 4496 790 4556
rect 830 4496 832 4556
rect 836 4496 840 4556
rect 844 4496 848 4556
rect 852 4498 854 4556
rect 931 4516 933 4556
rect 937 4516 943 4556
rect 947 4516 949 4556
rect 852 4496 866 4498
rect 1010 4496 1012 4556
rect 1016 4496 1020 4556
rect 1024 4496 1028 4556
rect 1032 4498 1034 4556
rect 1112 4516 1114 4556
rect 1118 4516 1122 4556
rect 1126 4516 1128 4556
rect 1140 4536 1144 4556
rect 1148 4536 1150 4556
rect 1032 4496 1046 4498
rect 1231 4516 1233 4556
rect 1237 4516 1243 4556
rect 1247 4516 1249 4556
rect 1303 4536 1305 4556
rect 1309 4536 1311 4556
rect 1323 4536 1325 4556
rect 1329 4536 1331 4556
rect 1383 4516 1385 4556
rect 1389 4516 1391 4556
rect 1403 4516 1405 4556
rect 1409 4528 1411 4556
rect 1423 4528 1425 4556
rect 1409 4516 1425 4528
rect 1429 4516 1431 4556
rect 1491 4516 1493 4556
rect 1497 4516 1503 4556
rect 1507 4516 1509 4556
rect 1549 4536 1551 4556
rect 1555 4536 1557 4556
rect 1569 4536 1571 4556
rect 1575 4536 1577 4556
rect 1630 4496 1632 4556
rect 1636 4496 1640 4556
rect 1644 4496 1648 4556
rect 1652 4498 1654 4556
rect 1750 4536 1752 4556
rect 1756 4536 1760 4556
rect 1652 4496 1666 4498
rect 1772 4516 1774 4556
rect 1778 4516 1782 4556
rect 1786 4516 1788 4556
rect 1829 4536 1831 4556
rect 1835 4536 1837 4556
rect 1903 4536 1905 4556
rect 1909 4536 1911 4556
rect 1952 4516 1954 4556
rect 1958 4516 1962 4556
rect 1966 4516 1968 4556
rect 1980 4536 1984 4556
rect 1988 4536 1990 4556
rect 2049 4536 2051 4556
rect 2055 4536 2057 4556
rect 2069 4536 2071 4556
rect 2075 4536 2077 4556
rect 2129 4536 2131 4556
rect 2135 4536 2137 4556
rect 2189 4516 2191 4556
rect 2195 4528 2197 4556
rect 2209 4528 2211 4556
rect 2195 4516 2211 4528
rect 2215 4516 2217 4556
rect 2229 4516 2231 4556
rect 2235 4516 2237 4556
rect 2303 4516 2305 4556
rect 2309 4544 2325 4556
rect 2309 4516 2311 4544
rect 2323 4516 2325 4544
rect 2329 4516 2331 4556
rect 2343 4516 2345 4556
rect 2349 4526 2351 4556
rect 2363 4526 2365 4556
rect 2349 4516 2365 4526
rect 2369 4516 2371 4556
rect 2409 4536 2411 4556
rect 2415 4536 2417 4556
rect 2429 4536 2431 4556
rect 2435 4536 2437 4556
rect 2449 4536 2451 4556
rect 2439 4516 2451 4536
rect 2455 4516 2457 4556
rect 2512 4516 2514 4556
rect 2518 4516 2522 4556
rect 2526 4516 2528 4556
rect 2540 4536 2544 4556
rect 2548 4536 2550 4556
rect 2644 4516 2646 4556
rect 2650 4516 2654 4556
rect 2658 4516 2660 4556
rect 2672 4516 2674 4556
rect 2678 4516 2682 4556
rect 2686 4516 2688 4556
rect 2733 4516 2735 4556
rect 2739 4536 2741 4556
rect 2753 4536 2755 4556
rect 2759 4536 2765 4556
rect 2769 4536 2773 4556
rect 2785 4536 2787 4556
rect 2791 4536 2797 4556
rect 2801 4536 2803 4556
rect 2815 4536 2819 4556
rect 2823 4536 2825 4556
rect 2863 4536 2865 4556
rect 2869 4536 2873 4556
rect 2877 4536 2879 4556
rect 2891 4536 2893 4556
rect 2897 4536 2903 4556
rect 2907 4536 2909 4556
rect 2921 4536 2925 4556
rect 2739 4516 2749 4536
rect 2912 4516 2925 4536
rect 2929 4516 2931 4556
rect 2983 4536 2985 4556
rect 2989 4536 2991 4556
rect 3043 4516 3045 4556
rect 3049 4516 3051 4556
rect 3063 4516 3065 4556
rect 3069 4528 3071 4556
rect 3083 4528 3085 4556
rect 3069 4516 3085 4528
rect 3089 4516 3091 4556
rect 3143 4536 3145 4556
rect 3149 4536 3151 4556
rect 3163 4536 3165 4556
rect 3169 4536 3171 4556
rect 3223 4516 3225 4556
rect 3229 4516 3231 4556
rect 3243 4516 3245 4556
rect 3249 4528 3251 4556
rect 3263 4528 3265 4556
rect 3249 4516 3265 4528
rect 3269 4516 3271 4556
rect 3323 4536 3325 4556
rect 3329 4536 3331 4556
rect 3343 4536 3345 4556
rect 3349 4536 3351 4556
rect 3403 4536 3405 4556
rect 3409 4536 3411 4556
rect 3449 4516 3451 4556
rect 3455 4536 3459 4556
rect 3471 4536 3473 4556
rect 3477 4536 3483 4556
rect 3487 4536 3489 4556
rect 3501 4536 3503 4556
rect 3507 4536 3511 4556
rect 3515 4536 3517 4556
rect 3555 4536 3557 4556
rect 3561 4536 3565 4556
rect 3577 4536 3579 4556
rect 3583 4536 3589 4556
rect 3593 4536 3595 4556
rect 3607 4536 3611 4556
rect 3615 4536 3621 4556
rect 3625 4536 3627 4556
rect 3639 4536 3641 4556
rect 3455 4516 3468 4536
rect 3631 4516 3641 4536
rect 3645 4516 3647 4556
rect 3689 4516 3691 4556
rect 3695 4528 3697 4556
rect 3709 4528 3711 4556
rect 3695 4516 3711 4528
rect 3715 4516 3717 4556
rect 3729 4516 3731 4556
rect 3735 4516 3737 4556
rect 3791 4516 3793 4556
rect 3797 4516 3803 4556
rect 3807 4516 3809 4556
rect 3883 4516 3885 4556
rect 3889 4516 3891 4556
rect 3903 4516 3905 4556
rect 3909 4516 3911 4556
rect 3923 4516 3925 4556
rect 3929 4516 3931 4556
rect 3943 4516 3945 4556
rect 3949 4516 3951 4556
rect 3963 4516 3965 4556
rect 3969 4516 3971 4556
rect 3983 4516 3985 4556
rect 3989 4516 3991 4556
rect 4003 4516 4005 4556
rect 4009 4516 4011 4556
rect 4023 4516 4025 4556
rect 4029 4516 4031 4556
rect 4081 4516 4083 4556
rect 4087 4516 4089 4556
rect 4101 4536 4105 4556
rect 4109 4536 4111 4556
rect 4151 4516 4153 4556
rect 4157 4516 4163 4556
rect 4167 4516 4169 4556
rect 4229 4536 4231 4556
rect 4235 4536 4237 4556
rect 4289 4516 4291 4556
rect 4295 4528 4297 4556
rect 4309 4528 4311 4556
rect 4295 4516 4311 4528
rect 4315 4516 4317 4556
rect 4329 4516 4331 4556
rect 4335 4516 4337 4556
rect 4389 4516 4391 4556
rect 4395 4536 4399 4556
rect 4411 4536 4413 4556
rect 4417 4536 4423 4556
rect 4427 4536 4429 4556
rect 4441 4536 4443 4556
rect 4447 4536 4451 4556
rect 4455 4536 4457 4556
rect 4495 4536 4497 4556
rect 4501 4536 4505 4556
rect 4517 4536 4519 4556
rect 4523 4536 4529 4556
rect 4533 4536 4535 4556
rect 4547 4536 4551 4556
rect 4555 4536 4561 4556
rect 4565 4536 4567 4556
rect 4579 4536 4581 4556
rect 4395 4516 4408 4536
rect 4571 4516 4581 4536
rect 4585 4516 4587 4556
rect 4629 4536 4631 4556
rect 4635 4536 4639 4556
rect 4651 4516 4653 4556
rect 4657 4516 4659 4556
rect 4711 4516 4713 4556
rect 4717 4516 4723 4556
rect 4727 4516 4729 4556
rect 51 4104 53 4144
rect 57 4104 63 4144
rect 67 4104 69 4144
rect 112 4104 114 4144
rect 118 4104 122 4144
rect 126 4104 128 4144
rect 140 4104 144 4124
rect 148 4104 150 4124
rect 231 4104 233 4144
rect 237 4104 243 4144
rect 247 4104 249 4144
rect 303 4104 305 4124
rect 309 4104 311 4124
rect 323 4104 325 4124
rect 329 4104 331 4124
rect 383 4104 385 4144
rect 389 4104 391 4144
rect 403 4104 405 4144
rect 409 4132 425 4144
rect 409 4104 411 4132
rect 423 4104 425 4132
rect 429 4104 431 4144
rect 469 4104 471 4144
rect 475 4132 491 4144
rect 475 4104 477 4132
rect 489 4104 491 4132
rect 495 4104 497 4144
rect 509 4104 511 4144
rect 515 4104 517 4144
rect 583 4104 585 4124
rect 589 4104 591 4124
rect 650 4104 652 4124
rect 656 4104 660 4124
rect 672 4104 674 4144
rect 678 4104 682 4144
rect 686 4104 688 4144
rect 743 4104 745 4124
rect 749 4104 751 4124
rect 790 4104 792 4164
rect 796 4104 800 4164
rect 804 4104 808 4164
rect 812 4162 826 4164
rect 812 4104 814 4162
rect 1034 4162 1048 4164
rect 924 4104 926 4144
rect 930 4104 934 4144
rect 938 4104 940 4144
rect 952 4104 954 4144
rect 958 4104 962 4144
rect 966 4104 968 4144
rect 1046 4104 1048 4162
rect 1052 4104 1056 4164
rect 1060 4104 1064 4164
rect 1068 4104 1070 4164
rect 1110 4104 1112 4164
rect 1116 4104 1120 4164
rect 1124 4104 1128 4164
rect 1132 4162 1146 4164
rect 1132 4104 1134 4162
rect 1314 4162 1328 4164
rect 1231 4104 1233 4144
rect 1237 4104 1243 4144
rect 1247 4104 1249 4144
rect 1326 4104 1328 4162
rect 1332 4104 1336 4164
rect 1340 4104 1344 4164
rect 1348 4104 1350 4164
rect 1411 4104 1413 4144
rect 1417 4104 1423 4144
rect 1427 4104 1429 4144
rect 1470 4104 1472 4164
rect 1476 4104 1480 4164
rect 1484 4104 1488 4164
rect 1492 4162 1506 4164
rect 1492 4104 1494 4162
rect 1583 4104 1585 4124
rect 1589 4104 1591 4124
rect 1603 4104 1605 4124
rect 1609 4104 1611 4124
rect 1663 4104 1665 4124
rect 1669 4104 1671 4124
rect 1683 4104 1685 4124
rect 1689 4104 1691 4124
rect 1729 4104 1731 4144
rect 1735 4132 1751 4144
rect 1735 4104 1737 4132
rect 1749 4104 1751 4132
rect 1755 4104 1757 4144
rect 1769 4104 1771 4144
rect 1775 4104 1777 4144
rect 1851 4104 1853 4144
rect 1857 4104 1863 4144
rect 1867 4104 1869 4144
rect 1909 4104 1911 4124
rect 1915 4104 1917 4124
rect 1970 4104 1972 4164
rect 1976 4104 1980 4164
rect 1984 4104 1988 4164
rect 1992 4162 2006 4164
rect 1992 4104 1994 4162
rect 2070 4104 2072 4164
rect 2076 4104 2080 4164
rect 2084 4104 2088 4164
rect 2092 4162 2106 4164
rect 2092 4104 2094 4162
rect 2173 4104 2175 4144
rect 2179 4124 2189 4144
rect 2352 4124 2365 4144
rect 2179 4104 2181 4124
rect 2193 4104 2195 4124
rect 2199 4104 2205 4124
rect 2209 4104 2213 4124
rect 2225 4104 2227 4124
rect 2231 4104 2237 4124
rect 2241 4104 2243 4124
rect 2255 4104 2259 4124
rect 2263 4104 2265 4124
rect 2303 4104 2305 4124
rect 2309 4104 2313 4124
rect 2317 4104 2319 4124
rect 2331 4104 2333 4124
rect 2337 4104 2343 4124
rect 2347 4104 2349 4124
rect 2361 4104 2365 4124
rect 2369 4104 2371 4144
rect 2409 4104 2411 4124
rect 2415 4104 2419 4124
rect 2431 4104 2433 4144
rect 2437 4104 2439 4144
rect 2503 4104 2505 4124
rect 2509 4104 2511 4124
rect 2563 4104 2565 4124
rect 2569 4104 2571 4124
rect 2583 4104 2585 4124
rect 2589 4104 2591 4124
rect 2629 4104 2631 4144
rect 2635 4124 2648 4144
rect 2811 4124 2821 4144
rect 2635 4104 2639 4124
rect 2651 4104 2653 4124
rect 2657 4104 2663 4124
rect 2667 4104 2669 4124
rect 2681 4104 2683 4124
rect 2687 4104 2691 4124
rect 2695 4104 2697 4124
rect 2735 4104 2737 4124
rect 2741 4104 2745 4124
rect 2757 4104 2759 4124
rect 2763 4104 2769 4124
rect 2773 4104 2775 4124
rect 2787 4104 2791 4124
rect 2795 4104 2801 4124
rect 2805 4104 2807 4124
rect 2819 4104 2821 4124
rect 2825 4104 2827 4144
rect 2869 4104 2871 4124
rect 2875 4104 2877 4124
rect 2943 4104 2945 4124
rect 2949 4104 2951 4124
rect 2963 4104 2965 4124
rect 2969 4104 2971 4124
rect 3009 4104 3011 4144
rect 3015 4132 3031 4144
rect 3015 4104 3017 4132
rect 3029 4104 3031 4132
rect 3035 4104 3037 4144
rect 3049 4104 3051 4144
rect 3055 4104 3057 4144
rect 3111 4104 3113 4144
rect 3117 4104 3123 4144
rect 3127 4104 3129 4144
rect 3211 4104 3213 4144
rect 3217 4104 3223 4144
rect 3227 4104 3229 4144
rect 3291 4104 3293 4144
rect 3297 4104 3303 4144
rect 3307 4104 3309 4144
rect 3349 4104 3351 4124
rect 3355 4104 3357 4124
rect 3369 4104 3371 4124
rect 3375 4104 3377 4124
rect 3433 4104 3435 4144
rect 3439 4124 3449 4144
rect 3612 4124 3625 4144
rect 3439 4104 3441 4124
rect 3453 4104 3455 4124
rect 3459 4104 3465 4124
rect 3469 4104 3473 4124
rect 3485 4104 3487 4124
rect 3491 4104 3497 4124
rect 3501 4104 3503 4124
rect 3515 4104 3519 4124
rect 3523 4104 3525 4124
rect 3563 4104 3565 4124
rect 3569 4104 3573 4124
rect 3577 4104 3579 4124
rect 3591 4104 3593 4124
rect 3597 4104 3603 4124
rect 3607 4104 3609 4124
rect 3621 4104 3625 4124
rect 3629 4104 3631 4144
rect 3691 4104 3693 4144
rect 3697 4104 3703 4144
rect 3707 4104 3709 4144
rect 3749 4104 3751 4124
rect 3755 4104 3757 4124
rect 3769 4104 3771 4124
rect 3775 4104 3777 4124
rect 3829 4104 3831 4144
rect 3835 4124 3848 4144
rect 4011 4124 4021 4144
rect 3835 4104 3839 4124
rect 3851 4104 3853 4124
rect 3857 4104 3863 4124
rect 3867 4104 3869 4124
rect 3881 4104 3883 4124
rect 3887 4104 3891 4124
rect 3895 4104 3897 4124
rect 3935 4104 3937 4124
rect 3941 4104 3945 4124
rect 3957 4104 3959 4124
rect 3963 4104 3969 4124
rect 3973 4104 3975 4124
rect 3987 4104 3991 4124
rect 3995 4104 4001 4124
rect 4005 4104 4007 4124
rect 4019 4104 4021 4124
rect 4025 4104 4027 4144
rect 4069 4104 4071 4124
rect 4075 4104 4077 4124
rect 4089 4104 4091 4124
rect 4095 4104 4097 4124
rect 4170 4104 4172 4124
rect 4176 4104 4180 4124
rect 4192 4104 4194 4144
rect 4198 4104 4202 4144
rect 4206 4104 4208 4144
rect 4249 4104 4251 4124
rect 4255 4104 4259 4124
rect 4271 4104 4273 4144
rect 4277 4104 4279 4144
rect 4343 4104 4345 4124
rect 4349 4104 4351 4124
rect 4363 4104 4365 4124
rect 4369 4104 4371 4124
rect 4430 4104 4432 4124
rect 4436 4104 4440 4124
rect 4452 4104 4454 4144
rect 4458 4104 4462 4144
rect 4466 4104 4468 4144
rect 4509 4104 4511 4144
rect 4515 4124 4528 4144
rect 4691 4124 4701 4144
rect 4515 4104 4519 4124
rect 4531 4104 4533 4124
rect 4537 4104 4543 4124
rect 4547 4104 4549 4124
rect 4561 4104 4563 4124
rect 4567 4104 4571 4124
rect 4575 4104 4577 4124
rect 4615 4104 4617 4124
rect 4621 4104 4625 4124
rect 4637 4104 4639 4124
rect 4643 4104 4649 4124
rect 4653 4104 4655 4124
rect 4667 4104 4671 4124
rect 4675 4104 4681 4124
rect 4685 4104 4687 4124
rect 4699 4104 4701 4124
rect 4705 4104 4707 4144
rect 51 4036 53 4076
rect 57 4036 63 4076
rect 67 4036 69 4076
rect 111 4036 113 4076
rect 117 4036 123 4076
rect 127 4036 129 4076
rect 211 4036 213 4076
rect 217 4036 223 4076
rect 227 4036 229 4076
rect 283 4036 285 4076
rect 289 4036 291 4076
rect 303 4036 305 4076
rect 309 4048 311 4076
rect 323 4048 325 4076
rect 309 4036 325 4048
rect 329 4036 331 4076
rect 372 4036 374 4076
rect 378 4036 382 4076
rect 386 4036 388 4076
rect 400 4056 404 4076
rect 408 4056 410 4076
rect 483 4056 485 4076
rect 489 4056 491 4076
rect 503 4056 505 4076
rect 509 4056 511 4076
rect 551 4036 553 4076
rect 557 4036 563 4076
rect 567 4036 569 4076
rect 629 4036 631 4076
rect 635 4048 637 4076
rect 649 4048 651 4076
rect 635 4036 651 4048
rect 655 4036 657 4076
rect 669 4036 671 4076
rect 675 4036 677 4076
rect 766 4018 768 4076
rect 754 4016 768 4018
rect 772 4016 776 4076
rect 780 4016 784 4076
rect 788 4016 790 4076
rect 830 4016 832 4076
rect 836 4016 840 4076
rect 844 4016 848 4076
rect 852 4018 854 4076
rect 943 4036 945 4076
rect 949 4036 951 4076
rect 963 4036 965 4076
rect 969 4048 971 4076
rect 983 4048 985 4076
rect 969 4036 985 4048
rect 989 4036 991 4076
rect 1029 4036 1031 4076
rect 1035 4048 1037 4076
rect 1049 4048 1051 4076
rect 1035 4036 1051 4048
rect 1055 4036 1057 4076
rect 1069 4036 1071 4076
rect 1075 4036 1077 4076
rect 1143 4056 1145 4076
rect 1149 4056 1151 4076
rect 852 4016 866 4018
rect 1226 4018 1228 4076
rect 1214 4016 1228 4018
rect 1232 4016 1236 4076
rect 1240 4016 1244 4076
rect 1248 4016 1250 4076
rect 1289 4056 1291 4076
rect 1295 4056 1297 4076
rect 1350 4016 1352 4076
rect 1356 4016 1360 4076
rect 1364 4016 1368 4076
rect 1372 4018 1374 4076
rect 1372 4016 1386 4018
rect 1450 4016 1452 4076
rect 1456 4016 1460 4076
rect 1464 4016 1468 4076
rect 1472 4018 1474 4076
rect 1551 4036 1553 4076
rect 1557 4036 1563 4076
rect 1567 4036 1569 4076
rect 1643 4056 1645 4076
rect 1649 4056 1651 4076
rect 1663 4056 1665 4076
rect 1669 4056 1671 4076
rect 1472 4016 1486 4018
rect 1733 4036 1735 4076
rect 1739 4036 1741 4076
rect 1753 4036 1755 4076
rect 1759 4036 1765 4076
rect 1769 4036 1771 4076
rect 1823 4036 1825 4076
rect 1829 4036 1831 4076
rect 1843 4036 1845 4076
rect 1849 4048 1851 4076
rect 1863 4048 1865 4076
rect 1849 4036 1865 4048
rect 1869 4036 1871 4076
rect 1909 4056 1911 4076
rect 1915 4056 1917 4076
rect 1929 4056 1931 4076
rect 1935 4056 1937 4076
rect 2003 4056 2005 4076
rect 2009 4056 2011 4076
rect 2049 4036 2051 4076
rect 2055 4048 2057 4076
rect 2069 4048 2071 4076
rect 2055 4036 2071 4048
rect 2075 4036 2077 4076
rect 2089 4036 2091 4076
rect 2095 4036 2097 4076
rect 2149 4056 2151 4076
rect 2155 4056 2157 4076
rect 2211 4036 2213 4076
rect 2217 4036 2223 4076
rect 2227 4036 2229 4076
rect 2290 4016 2292 4076
rect 2296 4016 2300 4076
rect 2304 4016 2308 4076
rect 2312 4018 2314 4076
rect 2389 4056 2391 4076
rect 2395 4056 2399 4076
rect 2312 4016 2326 4018
rect 2411 4036 2413 4076
rect 2417 4036 2419 4076
rect 2469 4036 2471 4076
rect 2475 4036 2477 4076
rect 2489 4036 2491 4076
rect 2495 4036 2497 4076
rect 2509 4036 2511 4076
rect 2515 4036 2517 4076
rect 2529 4036 2531 4076
rect 2535 4036 2537 4076
rect 2549 4036 2551 4076
rect 2555 4036 2557 4076
rect 2569 4036 2571 4076
rect 2575 4036 2577 4076
rect 2589 4036 2591 4076
rect 2595 4036 2597 4076
rect 2609 4036 2611 4076
rect 2615 4036 2617 4076
rect 2673 4036 2675 4076
rect 2679 4056 2681 4076
rect 2693 4056 2695 4076
rect 2699 4056 2705 4076
rect 2709 4056 2713 4076
rect 2725 4056 2727 4076
rect 2731 4056 2737 4076
rect 2741 4056 2743 4076
rect 2755 4056 2759 4076
rect 2763 4056 2765 4076
rect 2803 4056 2805 4076
rect 2809 4056 2813 4076
rect 2817 4056 2819 4076
rect 2831 4056 2833 4076
rect 2837 4056 2843 4076
rect 2847 4056 2849 4076
rect 2861 4056 2865 4076
rect 2679 4036 2689 4056
rect 2852 4036 2865 4056
rect 2869 4036 2871 4076
rect 2909 4056 2911 4076
rect 2915 4056 2917 4076
rect 2969 4036 2971 4076
rect 2975 4048 2977 4076
rect 2989 4048 2991 4076
rect 2975 4036 2991 4048
rect 2995 4036 2997 4076
rect 3009 4036 3011 4076
rect 3015 4036 3017 4076
rect 3069 4056 3071 4076
rect 3075 4056 3077 4076
rect 3089 4056 3091 4076
rect 3095 4056 3097 4076
rect 3151 4036 3153 4076
rect 3157 4036 3163 4076
rect 3167 4036 3169 4076
rect 3250 4056 3252 4076
rect 3256 4056 3260 4076
rect 3272 4036 3274 4076
rect 3278 4036 3282 4076
rect 3286 4036 3288 4076
rect 3329 4036 3331 4076
rect 3335 4036 3341 4076
rect 3345 4036 3347 4076
rect 3359 4036 3361 4076
rect 3365 4036 3367 4076
rect 3443 4056 3445 4076
rect 3449 4056 3451 4076
rect 3463 4056 3465 4076
rect 3469 4056 3471 4076
rect 3523 4056 3525 4076
rect 3529 4056 3531 4076
rect 3569 4036 3571 4076
rect 3575 4056 3579 4076
rect 3591 4056 3593 4076
rect 3597 4056 3603 4076
rect 3607 4056 3609 4076
rect 3621 4056 3623 4076
rect 3627 4056 3631 4076
rect 3635 4056 3637 4076
rect 3675 4056 3677 4076
rect 3681 4056 3685 4076
rect 3697 4056 3699 4076
rect 3703 4056 3709 4076
rect 3713 4056 3715 4076
rect 3727 4056 3731 4076
rect 3735 4056 3741 4076
rect 3745 4056 3747 4076
rect 3759 4056 3761 4076
rect 3575 4036 3588 4056
rect 3751 4036 3761 4056
rect 3765 4036 3767 4076
rect 3830 4056 3832 4076
rect 3836 4056 3840 4076
rect 3852 4036 3854 4076
rect 3858 4036 3862 4076
rect 3866 4036 3868 4076
rect 3909 4056 3911 4076
rect 3915 4056 3917 4076
rect 3929 4056 3931 4076
rect 3935 4056 3937 4076
rect 4003 4056 4005 4076
rect 4009 4056 4011 4076
rect 4023 4056 4025 4076
rect 4029 4056 4031 4076
rect 4069 4036 4071 4076
rect 4075 4036 4081 4076
rect 4085 4036 4087 4076
rect 4099 4036 4101 4076
rect 4105 4036 4107 4076
rect 4169 4036 4171 4076
rect 4175 4048 4177 4076
rect 4189 4048 4191 4076
rect 4175 4036 4191 4048
rect 4195 4036 4197 4076
rect 4209 4036 4211 4076
rect 4215 4036 4217 4076
rect 4283 4036 4285 4076
rect 4289 4036 4291 4076
rect 4303 4036 4305 4076
rect 4309 4048 4311 4076
rect 4323 4048 4325 4076
rect 4309 4036 4325 4048
rect 4329 4036 4331 4076
rect 4383 4056 4385 4076
rect 4389 4056 4391 4076
rect 4429 4036 4431 4076
rect 4435 4056 4439 4076
rect 4451 4056 4453 4076
rect 4457 4056 4463 4076
rect 4467 4056 4469 4076
rect 4481 4056 4483 4076
rect 4487 4056 4491 4076
rect 4495 4056 4497 4076
rect 4535 4056 4537 4076
rect 4541 4056 4545 4076
rect 4557 4056 4559 4076
rect 4563 4056 4569 4076
rect 4573 4056 4575 4076
rect 4587 4056 4591 4076
rect 4595 4056 4601 4076
rect 4605 4056 4607 4076
rect 4619 4056 4621 4076
rect 4435 4036 4448 4056
rect 4611 4036 4621 4056
rect 4625 4036 4627 4076
rect 4669 4056 4671 4076
rect 4675 4056 4677 4076
rect 43 3624 45 3644
rect 49 3624 51 3644
rect 63 3624 65 3644
rect 69 3624 71 3644
rect 109 3624 111 3664
rect 115 3652 131 3664
rect 115 3624 117 3652
rect 129 3624 131 3652
rect 135 3624 137 3664
rect 149 3624 151 3664
rect 155 3624 157 3664
rect 223 3624 225 3644
rect 229 3624 231 3644
rect 290 3624 292 3644
rect 296 3624 300 3644
rect 312 3624 314 3664
rect 318 3624 322 3664
rect 326 3624 328 3664
rect 393 3624 395 3664
rect 399 3624 401 3664
rect 413 3624 415 3664
rect 419 3624 425 3664
rect 429 3624 431 3664
rect 491 3624 493 3664
rect 497 3624 503 3664
rect 507 3624 509 3664
rect 571 3624 573 3664
rect 577 3624 583 3664
rect 587 3624 589 3664
rect 894 3682 908 3684
rect 629 3624 631 3644
rect 635 3624 637 3644
rect 689 3624 691 3664
rect 695 3652 711 3664
rect 695 3624 697 3652
rect 709 3624 711 3652
rect 715 3624 717 3664
rect 729 3624 731 3664
rect 735 3624 737 3664
rect 791 3624 793 3664
rect 797 3624 803 3664
rect 807 3624 809 3664
rect 906 3624 908 3682
rect 912 3624 916 3684
rect 920 3624 924 3684
rect 928 3624 930 3684
rect 972 3624 974 3664
rect 978 3624 982 3664
rect 986 3624 988 3664
rect 1000 3624 1004 3644
rect 1008 3624 1010 3644
rect 1070 3624 1072 3684
rect 1076 3624 1080 3684
rect 1084 3624 1088 3684
rect 1092 3682 1106 3684
rect 1092 3624 1094 3682
rect 1172 3624 1174 3664
rect 1178 3624 1182 3664
rect 1186 3624 1188 3664
rect 1354 3682 1368 3684
rect 1200 3624 1204 3644
rect 1208 3624 1210 3644
rect 1269 3624 1271 3644
rect 1275 3624 1277 3644
rect 1366 3624 1368 3682
rect 1372 3624 1376 3684
rect 1380 3624 1384 3684
rect 1388 3624 1390 3684
rect 1443 3624 1445 3644
rect 1449 3624 1451 3644
rect 1503 3624 1505 3664
rect 1509 3624 1511 3664
rect 1523 3624 1525 3664
rect 1529 3652 1545 3664
rect 1529 3624 1531 3652
rect 1543 3624 1545 3652
rect 1549 3624 1551 3664
rect 1603 3624 1605 3644
rect 1609 3624 1611 3644
rect 1652 3624 1654 3664
rect 1658 3624 1662 3664
rect 1666 3624 1668 3664
rect 1680 3624 1684 3644
rect 1688 3624 1690 3644
rect 1749 3624 1751 3644
rect 1755 3624 1757 3644
rect 1769 3624 1771 3644
rect 1775 3624 1777 3644
rect 1850 3624 1852 3644
rect 1856 3624 1860 3644
rect 1872 3624 1874 3664
rect 1878 3624 1882 3664
rect 1886 3624 1888 3664
rect 1951 3624 1953 3664
rect 1957 3624 1963 3664
rect 1967 3624 1969 3664
rect 2039 3644 2051 3664
rect 2009 3624 2011 3644
rect 2015 3624 2017 3644
rect 2029 3624 2031 3644
rect 2035 3624 2037 3644
rect 2049 3624 2051 3644
rect 2055 3624 2057 3664
rect 2109 3624 2111 3644
rect 2115 3624 2119 3644
rect 2131 3624 2133 3664
rect 2137 3624 2139 3664
rect 2203 3624 2205 3664
rect 2209 3624 2211 3664
rect 2223 3624 2225 3664
rect 2229 3624 2231 3664
rect 2243 3624 2245 3664
rect 2249 3624 2251 3664
rect 2263 3624 2265 3664
rect 2269 3624 2271 3664
rect 2283 3624 2285 3664
rect 2289 3624 2291 3664
rect 2303 3624 2305 3664
rect 2309 3624 2311 3664
rect 2323 3624 2325 3664
rect 2329 3624 2331 3664
rect 2343 3624 2345 3664
rect 2349 3624 2351 3664
rect 2393 3624 2395 3664
rect 2399 3644 2409 3664
rect 2572 3644 2585 3664
rect 2399 3624 2401 3644
rect 2413 3624 2415 3644
rect 2419 3624 2425 3644
rect 2429 3624 2433 3644
rect 2445 3624 2447 3644
rect 2451 3624 2457 3644
rect 2461 3624 2463 3644
rect 2475 3624 2479 3644
rect 2483 3624 2485 3644
rect 2523 3624 2525 3644
rect 2529 3624 2533 3644
rect 2537 3624 2539 3644
rect 2551 3624 2553 3644
rect 2557 3624 2563 3644
rect 2567 3624 2569 3644
rect 2581 3624 2585 3644
rect 2589 3624 2591 3664
rect 2643 3624 2645 3664
rect 2649 3624 2651 3664
rect 2663 3624 2665 3664
rect 2669 3652 2685 3664
rect 2669 3624 2671 3652
rect 2683 3624 2685 3652
rect 2689 3624 2691 3664
rect 2743 3624 2745 3644
rect 2749 3624 2751 3644
rect 2803 3624 2805 3644
rect 2809 3624 2811 3644
rect 2823 3624 2825 3644
rect 2829 3624 2831 3644
rect 2883 3624 2885 3644
rect 2889 3624 2891 3644
rect 2903 3624 2905 3644
rect 2909 3624 2911 3644
rect 2963 3624 2965 3644
rect 2969 3624 2971 3644
rect 2983 3624 2985 3644
rect 2989 3624 2991 3644
rect 3029 3624 3031 3644
rect 3035 3624 3037 3644
rect 3103 3624 3105 3644
rect 3109 3624 3111 3644
rect 3149 3624 3151 3664
rect 3155 3652 3171 3664
rect 3155 3624 3157 3652
rect 3169 3624 3171 3652
rect 3175 3624 3177 3664
rect 3189 3624 3191 3664
rect 3195 3624 3197 3664
rect 3270 3624 3272 3644
rect 3276 3624 3280 3644
rect 3292 3624 3294 3664
rect 3298 3624 3302 3664
rect 3306 3624 3308 3664
rect 3352 3624 3354 3664
rect 3358 3624 3362 3664
rect 3366 3624 3368 3664
rect 3380 3624 3384 3644
rect 3388 3624 3390 3644
rect 3449 3624 3451 3644
rect 3455 3624 3457 3644
rect 3509 3624 3511 3664
rect 3515 3624 3521 3664
rect 3525 3624 3527 3664
rect 3539 3624 3541 3664
rect 3545 3624 3547 3664
rect 3609 3624 3611 3664
rect 3615 3652 3631 3664
rect 3615 3624 3617 3652
rect 3629 3624 3631 3652
rect 3635 3624 3637 3664
rect 3649 3624 3651 3664
rect 3655 3624 3657 3664
rect 3709 3624 3711 3664
rect 3715 3652 3731 3664
rect 3715 3624 3717 3652
rect 3729 3624 3731 3652
rect 3735 3624 3737 3664
rect 3749 3624 3751 3664
rect 3755 3624 3757 3664
rect 3813 3624 3815 3664
rect 3819 3644 3829 3664
rect 3992 3644 4005 3664
rect 3819 3624 3821 3644
rect 3833 3624 3835 3644
rect 3839 3624 3845 3644
rect 3849 3624 3853 3644
rect 3865 3624 3867 3644
rect 3871 3624 3877 3644
rect 3881 3624 3883 3644
rect 3895 3624 3899 3644
rect 3903 3624 3905 3644
rect 3943 3624 3945 3644
rect 3949 3624 3953 3644
rect 3957 3624 3959 3644
rect 3971 3624 3973 3644
rect 3977 3624 3983 3644
rect 3987 3624 3989 3644
rect 4001 3624 4005 3644
rect 4009 3624 4011 3664
rect 4049 3624 4051 3644
rect 4055 3624 4059 3644
rect 4071 3624 4073 3664
rect 4077 3624 4079 3664
rect 4143 3624 4145 3644
rect 4149 3624 4151 3644
rect 4163 3624 4165 3644
rect 4169 3624 4171 3644
rect 4212 3624 4214 3664
rect 4218 3624 4222 3664
rect 4226 3624 4228 3664
rect 4240 3624 4244 3644
rect 4248 3624 4250 3644
rect 4309 3624 4311 3664
rect 4315 3644 4328 3664
rect 4491 3644 4501 3664
rect 4315 3624 4319 3644
rect 4331 3624 4333 3644
rect 4337 3624 4343 3644
rect 4347 3624 4349 3644
rect 4361 3624 4363 3644
rect 4367 3624 4371 3644
rect 4375 3624 4377 3644
rect 4415 3624 4417 3644
rect 4421 3624 4425 3644
rect 4437 3624 4439 3644
rect 4443 3624 4449 3644
rect 4453 3624 4455 3644
rect 4467 3624 4471 3644
rect 4475 3624 4481 3644
rect 4485 3624 4487 3644
rect 4499 3624 4501 3644
rect 4505 3624 4507 3664
rect 4549 3624 4551 3644
rect 4555 3624 4559 3644
rect 4571 3624 4573 3664
rect 4577 3624 4579 3664
rect 4643 3624 4645 3644
rect 4649 3624 4651 3644
rect 4689 3624 4691 3644
rect 4695 3624 4697 3644
rect 51 3556 53 3596
rect 57 3556 63 3596
rect 67 3556 69 3596
rect 113 3556 115 3596
rect 119 3576 121 3596
rect 133 3576 135 3596
rect 139 3576 145 3596
rect 149 3576 153 3596
rect 165 3576 167 3596
rect 171 3576 177 3596
rect 181 3576 183 3596
rect 195 3576 199 3596
rect 203 3576 205 3596
rect 243 3576 245 3596
rect 249 3576 253 3596
rect 257 3576 259 3596
rect 271 3576 273 3596
rect 277 3576 283 3596
rect 287 3576 289 3596
rect 301 3576 305 3596
rect 119 3556 129 3576
rect 292 3556 305 3576
rect 309 3556 311 3596
rect 363 3576 365 3596
rect 369 3576 371 3596
rect 431 3556 433 3596
rect 437 3556 443 3596
rect 447 3556 449 3596
rect 503 3556 505 3596
rect 509 3556 511 3596
rect 523 3556 525 3596
rect 529 3568 531 3596
rect 543 3568 545 3596
rect 529 3556 545 3568
rect 549 3556 551 3596
rect 603 3556 605 3596
rect 609 3556 611 3596
rect 623 3556 625 3596
rect 629 3568 631 3596
rect 643 3568 645 3596
rect 629 3556 645 3568
rect 649 3556 651 3596
rect 691 3556 693 3596
rect 697 3556 703 3596
rect 707 3556 709 3596
rect 769 3556 771 3596
rect 775 3566 777 3596
rect 789 3566 791 3596
rect 775 3556 791 3566
rect 795 3556 797 3596
rect 809 3556 811 3596
rect 815 3584 831 3596
rect 815 3556 817 3584
rect 829 3556 831 3584
rect 835 3556 837 3596
rect 889 3576 891 3596
rect 895 3576 897 3596
rect 986 3538 988 3596
rect 974 3536 988 3538
rect 992 3536 996 3596
rect 1000 3536 1004 3596
rect 1008 3536 1010 3596
rect 1052 3556 1054 3596
rect 1058 3556 1062 3596
rect 1066 3556 1068 3596
rect 1080 3576 1084 3596
rect 1088 3576 1090 3596
rect 1149 3576 1151 3596
rect 1155 3576 1157 3596
rect 1169 3576 1171 3596
rect 1175 3576 1177 3596
rect 1231 3556 1233 3596
rect 1237 3556 1243 3596
rect 1247 3556 1249 3596
rect 1311 3556 1313 3596
rect 1317 3556 1323 3596
rect 1327 3556 1329 3596
rect 1389 3556 1391 3596
rect 1395 3568 1397 3596
rect 1409 3568 1411 3596
rect 1395 3556 1411 3568
rect 1415 3556 1417 3596
rect 1429 3556 1431 3596
rect 1435 3556 1437 3596
rect 1493 3556 1495 3596
rect 1499 3576 1501 3596
rect 1513 3576 1515 3596
rect 1519 3576 1525 3596
rect 1529 3576 1533 3596
rect 1545 3576 1547 3596
rect 1551 3576 1557 3596
rect 1561 3576 1563 3596
rect 1575 3576 1579 3596
rect 1583 3576 1585 3596
rect 1623 3576 1625 3596
rect 1629 3576 1633 3596
rect 1637 3576 1639 3596
rect 1651 3576 1653 3596
rect 1657 3576 1663 3596
rect 1667 3576 1669 3596
rect 1681 3576 1685 3596
rect 1499 3556 1509 3576
rect 1672 3556 1685 3576
rect 1689 3556 1691 3596
rect 1751 3556 1753 3596
rect 1757 3556 1763 3596
rect 1767 3556 1769 3596
rect 1809 3556 1811 3596
rect 1815 3568 1817 3596
rect 1829 3568 1831 3596
rect 1815 3556 1831 3568
rect 1835 3556 1837 3596
rect 1849 3556 1851 3596
rect 1855 3556 1857 3596
rect 1909 3556 1911 3596
rect 1915 3556 1917 3596
rect 1991 3556 1993 3596
rect 1997 3556 2003 3596
rect 2007 3556 2009 3596
rect 2073 3556 2075 3596
rect 2079 3556 2081 3596
rect 2093 3556 2095 3596
rect 2099 3556 2105 3596
rect 2109 3556 2111 3596
rect 2151 3556 2153 3596
rect 2157 3556 2163 3596
rect 2167 3556 2169 3596
rect 2230 3536 2232 3596
rect 2236 3536 2240 3596
rect 2244 3536 2248 3596
rect 2252 3538 2254 3596
rect 2329 3576 2331 3596
rect 2335 3576 2337 3596
rect 2389 3576 2391 3596
rect 2395 3576 2397 3596
rect 2252 3536 2266 3538
rect 2449 3556 2451 3596
rect 2455 3576 2459 3596
rect 2471 3576 2473 3596
rect 2477 3576 2483 3596
rect 2487 3576 2489 3596
rect 2501 3576 2503 3596
rect 2507 3576 2511 3596
rect 2515 3576 2517 3596
rect 2555 3576 2557 3596
rect 2561 3576 2565 3596
rect 2577 3576 2579 3596
rect 2583 3576 2589 3596
rect 2593 3576 2595 3596
rect 2607 3576 2611 3596
rect 2615 3576 2621 3596
rect 2625 3576 2627 3596
rect 2639 3576 2641 3596
rect 2455 3556 2468 3576
rect 2631 3556 2641 3576
rect 2645 3556 2647 3596
rect 2689 3556 2691 3596
rect 2695 3568 2697 3596
rect 2709 3568 2711 3596
rect 2695 3556 2711 3568
rect 2715 3556 2717 3596
rect 2729 3556 2731 3596
rect 2735 3556 2737 3596
rect 2789 3576 2791 3596
rect 2795 3576 2799 3596
rect 2811 3556 2813 3596
rect 2817 3556 2819 3596
rect 2871 3556 2873 3596
rect 2877 3556 2883 3596
rect 2887 3556 2889 3596
rect 2949 3556 2951 3596
rect 2955 3576 2959 3596
rect 2971 3576 2973 3596
rect 2977 3576 2983 3596
rect 2987 3576 2989 3596
rect 3001 3576 3003 3596
rect 3007 3576 3011 3596
rect 3015 3576 3017 3596
rect 3055 3576 3057 3596
rect 3061 3576 3065 3596
rect 3077 3576 3079 3596
rect 3083 3576 3089 3596
rect 3093 3576 3095 3596
rect 3107 3576 3111 3596
rect 3115 3576 3121 3596
rect 3125 3576 3127 3596
rect 3139 3576 3141 3596
rect 2955 3556 2968 3576
rect 3131 3556 3141 3576
rect 3145 3556 3147 3596
rect 3203 3556 3205 3596
rect 3209 3556 3211 3596
rect 3223 3556 3225 3596
rect 3229 3568 3231 3596
rect 3243 3568 3245 3596
rect 3229 3556 3245 3568
rect 3249 3556 3251 3596
rect 3303 3576 3305 3596
rect 3309 3576 3311 3596
rect 3349 3576 3351 3596
rect 3355 3576 3357 3596
rect 3369 3576 3371 3596
rect 3375 3576 3377 3596
rect 3429 3576 3431 3596
rect 3435 3576 3437 3596
rect 3503 3576 3505 3596
rect 3509 3576 3511 3596
rect 3523 3576 3525 3596
rect 3529 3576 3531 3596
rect 3572 3556 3574 3596
rect 3578 3556 3582 3596
rect 3586 3556 3588 3596
rect 3600 3576 3604 3596
rect 3608 3576 3610 3596
rect 3669 3576 3671 3596
rect 3675 3576 3677 3596
rect 3689 3576 3691 3596
rect 3695 3576 3697 3596
rect 3709 3576 3711 3596
rect 3699 3556 3711 3576
rect 3715 3556 3717 3596
rect 3804 3556 3806 3596
rect 3810 3556 3814 3596
rect 3818 3556 3820 3596
rect 3832 3556 3834 3596
rect 3838 3556 3842 3596
rect 3846 3556 3848 3596
rect 3911 3556 3913 3596
rect 3917 3556 3923 3596
rect 3927 3556 3929 3596
rect 3969 3556 3971 3596
rect 3975 3576 3979 3596
rect 3991 3576 3993 3596
rect 3997 3576 4003 3596
rect 4007 3576 4009 3596
rect 4021 3576 4023 3596
rect 4027 3576 4031 3596
rect 4035 3576 4037 3596
rect 4075 3576 4077 3596
rect 4081 3576 4085 3596
rect 4097 3576 4099 3596
rect 4103 3576 4109 3596
rect 4113 3576 4115 3596
rect 4127 3576 4131 3596
rect 4135 3576 4141 3596
rect 4145 3576 4147 3596
rect 4159 3576 4161 3596
rect 3975 3556 3988 3576
rect 4151 3556 4161 3576
rect 4165 3556 4167 3596
rect 4209 3556 4211 3596
rect 4215 3576 4219 3596
rect 4231 3576 4233 3596
rect 4237 3576 4243 3596
rect 4247 3576 4249 3596
rect 4261 3576 4263 3596
rect 4267 3576 4271 3596
rect 4275 3576 4277 3596
rect 4315 3576 4317 3596
rect 4321 3576 4325 3596
rect 4337 3576 4339 3596
rect 4343 3576 4349 3596
rect 4353 3576 4355 3596
rect 4367 3576 4371 3596
rect 4375 3576 4381 3596
rect 4385 3576 4387 3596
rect 4399 3576 4401 3596
rect 4215 3556 4228 3576
rect 4391 3556 4401 3576
rect 4405 3556 4407 3596
rect 4463 3556 4465 3596
rect 4469 3556 4471 3596
rect 4483 3556 4485 3596
rect 4489 3556 4491 3596
rect 4503 3556 4505 3596
rect 4509 3556 4511 3596
rect 4523 3556 4525 3596
rect 4529 3556 4531 3596
rect 4543 3556 4545 3596
rect 4549 3556 4551 3596
rect 4563 3556 4565 3596
rect 4569 3556 4571 3596
rect 4583 3556 4585 3596
rect 4589 3556 4591 3596
rect 4603 3556 4605 3596
rect 4609 3556 4611 3596
rect 4649 3556 4651 3596
rect 4655 3568 4657 3596
rect 4669 3568 4671 3596
rect 4655 3556 4671 3568
rect 4675 3556 4677 3596
rect 4689 3556 4691 3596
rect 4695 3556 4697 3596
rect 33 3144 35 3184
rect 39 3164 49 3184
rect 212 3164 225 3184
rect 39 3144 41 3164
rect 53 3144 55 3164
rect 59 3144 65 3164
rect 69 3144 73 3164
rect 85 3144 87 3164
rect 91 3144 97 3164
rect 101 3144 103 3164
rect 115 3144 119 3164
rect 123 3144 125 3164
rect 163 3144 165 3164
rect 169 3144 173 3164
rect 177 3144 179 3164
rect 191 3144 193 3164
rect 197 3144 203 3164
rect 207 3144 209 3164
rect 221 3144 225 3164
rect 229 3144 231 3184
rect 304 3144 306 3184
rect 310 3144 314 3184
rect 318 3144 320 3184
rect 332 3144 334 3184
rect 338 3144 342 3184
rect 346 3144 348 3184
rect 411 3144 413 3184
rect 417 3144 423 3184
rect 427 3144 429 3184
rect 469 3144 471 3184
rect 475 3164 488 3184
rect 1034 3202 1048 3204
rect 651 3164 661 3184
rect 475 3144 479 3164
rect 491 3144 493 3164
rect 497 3144 503 3164
rect 507 3144 509 3164
rect 521 3144 523 3164
rect 527 3144 531 3164
rect 535 3144 537 3164
rect 575 3144 577 3164
rect 581 3144 585 3164
rect 597 3144 599 3164
rect 603 3144 609 3164
rect 613 3144 615 3164
rect 627 3144 631 3164
rect 635 3144 641 3164
rect 645 3144 647 3164
rect 659 3144 661 3164
rect 665 3144 667 3184
rect 723 3144 725 3184
rect 729 3144 731 3184
rect 743 3144 745 3184
rect 749 3172 765 3184
rect 749 3144 751 3172
rect 763 3144 765 3172
rect 769 3144 771 3184
rect 844 3144 846 3184
rect 850 3144 854 3184
rect 858 3144 860 3184
rect 872 3144 874 3184
rect 878 3144 882 3184
rect 886 3144 888 3184
rect 931 3144 933 3184
rect 937 3144 943 3184
rect 947 3144 949 3184
rect 1046 3144 1048 3202
rect 1052 3144 1056 3204
rect 1060 3144 1064 3204
rect 1068 3144 1070 3204
rect 1133 3144 1135 3184
rect 1139 3144 1141 3184
rect 1153 3144 1155 3184
rect 1159 3144 1165 3184
rect 1169 3144 1171 3184
rect 1210 3144 1212 3204
rect 1216 3144 1220 3204
rect 1224 3144 1228 3204
rect 1232 3202 1246 3204
rect 1232 3144 1234 3202
rect 1309 3144 1311 3184
rect 1315 3172 1331 3184
rect 1315 3144 1317 3172
rect 1329 3144 1331 3172
rect 1335 3144 1337 3184
rect 1349 3144 1351 3184
rect 1355 3144 1357 3184
rect 1411 3144 1413 3184
rect 1417 3144 1423 3184
rect 1427 3144 1429 3184
rect 1503 3144 1505 3184
rect 1509 3164 1521 3184
rect 1509 3144 1511 3164
rect 1523 3144 1525 3164
rect 1529 3144 1531 3164
rect 1543 3144 1545 3164
rect 1549 3144 1551 3164
rect 1611 3144 1613 3184
rect 1617 3144 1623 3184
rect 1627 3144 1629 3184
rect 1669 3144 1671 3184
rect 1675 3172 1691 3184
rect 1675 3144 1677 3172
rect 1689 3144 1691 3172
rect 1695 3144 1697 3184
rect 1709 3144 1711 3184
rect 1715 3144 1717 3184
rect 1783 3144 1785 3184
rect 1789 3144 1791 3184
rect 1803 3144 1805 3184
rect 1809 3172 1825 3184
rect 1809 3144 1811 3172
rect 1823 3144 1825 3172
rect 1829 3144 1831 3184
rect 1871 3144 1873 3184
rect 1877 3144 1883 3184
rect 1887 3144 1889 3184
rect 1949 3144 1951 3184
rect 1955 3172 1971 3184
rect 1955 3144 1957 3172
rect 1969 3144 1971 3172
rect 1975 3144 1977 3184
rect 1989 3144 1991 3184
rect 1995 3144 1997 3184
rect 2063 3144 2065 3184
rect 2069 3144 2071 3184
rect 2083 3144 2085 3184
rect 2089 3172 2105 3184
rect 2089 3144 2091 3172
rect 2103 3144 2105 3172
rect 2109 3144 2111 3184
rect 2149 3144 2151 3164
rect 2155 3144 2157 3164
rect 2209 3144 2211 3184
rect 2215 3172 2231 3184
rect 2215 3144 2217 3172
rect 2229 3144 2231 3172
rect 2235 3144 2237 3184
rect 2249 3144 2251 3184
rect 2255 3144 2257 3184
rect 2323 3144 2325 3164
rect 2329 3144 2331 3164
rect 2371 3144 2373 3184
rect 2377 3144 2383 3184
rect 2387 3144 2389 3184
rect 2449 3144 2451 3184
rect 2455 3164 2468 3184
rect 2631 3164 2641 3184
rect 2455 3144 2459 3164
rect 2471 3144 2473 3164
rect 2477 3144 2483 3164
rect 2487 3144 2489 3164
rect 2501 3144 2503 3164
rect 2507 3144 2511 3164
rect 2515 3144 2517 3164
rect 2555 3144 2557 3164
rect 2561 3144 2565 3164
rect 2577 3144 2579 3164
rect 2583 3144 2589 3164
rect 2593 3144 2595 3164
rect 2607 3144 2611 3164
rect 2615 3144 2621 3164
rect 2625 3144 2627 3164
rect 2639 3144 2641 3164
rect 2645 3144 2647 3184
rect 2689 3144 2691 3164
rect 2695 3144 2699 3164
rect 2711 3144 2713 3184
rect 2717 3144 2719 3184
rect 2769 3144 2771 3184
rect 2775 3164 2788 3184
rect 2951 3164 2961 3184
rect 2775 3144 2779 3164
rect 2791 3144 2793 3164
rect 2797 3144 2803 3164
rect 2807 3144 2809 3164
rect 2821 3144 2823 3164
rect 2827 3144 2831 3164
rect 2835 3144 2837 3164
rect 2875 3144 2877 3164
rect 2881 3144 2885 3164
rect 2897 3144 2899 3164
rect 2903 3144 2909 3164
rect 2913 3144 2915 3164
rect 2927 3144 2931 3164
rect 2935 3144 2941 3164
rect 2945 3144 2947 3164
rect 2959 3144 2961 3164
rect 2965 3144 2967 3184
rect 3023 3144 3025 3184
rect 3029 3144 3031 3184
rect 3043 3144 3045 3184
rect 3049 3172 3065 3184
rect 3049 3144 3051 3172
rect 3063 3144 3065 3172
rect 3069 3144 3071 3184
rect 3123 3144 3125 3184
rect 3129 3144 3131 3184
rect 3143 3144 3145 3184
rect 3149 3172 3165 3184
rect 3149 3144 3151 3172
rect 3163 3144 3165 3172
rect 3169 3144 3171 3184
rect 3209 3144 3211 3184
rect 3215 3172 3231 3184
rect 3215 3144 3217 3172
rect 3229 3144 3231 3172
rect 3235 3144 3237 3184
rect 3249 3144 3251 3184
rect 3255 3144 3257 3184
rect 3323 3144 3325 3184
rect 3329 3144 3331 3184
rect 3343 3144 3345 3184
rect 3349 3172 3365 3184
rect 3349 3144 3351 3172
rect 3363 3144 3365 3172
rect 3369 3144 3371 3184
rect 3409 3144 3411 3184
rect 3415 3172 3431 3184
rect 3415 3144 3417 3172
rect 3429 3144 3431 3172
rect 3435 3144 3437 3184
rect 3449 3144 3451 3184
rect 3455 3144 3457 3184
rect 3511 3144 3513 3184
rect 3517 3144 3523 3184
rect 3527 3144 3529 3184
rect 3591 3144 3593 3184
rect 3597 3144 3603 3184
rect 3607 3144 3609 3184
rect 3671 3144 3673 3184
rect 3677 3144 3683 3184
rect 3687 3144 3689 3184
rect 3751 3144 3753 3184
rect 3757 3144 3763 3184
rect 3767 3144 3769 3184
rect 3829 3144 3831 3164
rect 3835 3144 3839 3164
rect 3851 3144 3853 3184
rect 3857 3144 3859 3184
rect 3931 3144 3933 3184
rect 3937 3144 3943 3184
rect 3947 3144 3949 3184
rect 4003 3144 4005 3164
rect 4009 3144 4011 3164
rect 4023 3144 4025 3164
rect 4029 3144 4031 3164
rect 4069 3144 4071 3164
rect 4075 3144 4079 3164
rect 4091 3144 4093 3184
rect 4097 3144 4099 3184
rect 4163 3144 4165 3164
rect 4169 3144 4171 3164
rect 4223 3144 4225 3184
rect 4229 3144 4231 3184
rect 4243 3144 4245 3184
rect 4249 3172 4265 3184
rect 4249 3144 4251 3172
rect 4263 3144 4265 3172
rect 4269 3144 4271 3184
rect 4323 3144 4325 3164
rect 4329 3144 4331 3164
rect 4369 3144 4371 3184
rect 4375 3172 4391 3184
rect 4375 3144 4377 3172
rect 4389 3144 4391 3172
rect 4395 3144 4397 3184
rect 4409 3144 4411 3184
rect 4415 3144 4417 3184
rect 4491 3144 4493 3184
rect 4497 3144 4503 3184
rect 4507 3144 4509 3184
rect 4553 3144 4555 3184
rect 4559 3164 4569 3184
rect 4732 3164 4745 3184
rect 4559 3144 4561 3164
rect 4573 3144 4575 3164
rect 4579 3144 4585 3164
rect 4589 3144 4593 3164
rect 4605 3144 4607 3164
rect 4611 3144 4617 3164
rect 4621 3144 4623 3164
rect 4635 3144 4639 3164
rect 4643 3144 4645 3164
rect 4683 3144 4685 3164
rect 4689 3144 4693 3164
rect 4697 3144 4699 3164
rect 4711 3144 4713 3164
rect 4717 3144 4723 3164
rect 4727 3144 4729 3164
rect 4741 3144 4745 3164
rect 4749 3144 4751 3184
rect 64 3076 66 3116
rect 70 3076 74 3116
rect 78 3076 80 3116
rect 92 3076 94 3116
rect 98 3076 102 3116
rect 106 3076 108 3116
rect 173 3076 175 3116
rect 179 3076 181 3116
rect 193 3076 195 3116
rect 199 3076 205 3116
rect 209 3076 211 3116
rect 249 3076 251 3116
rect 255 3096 259 3116
rect 271 3096 273 3116
rect 277 3096 283 3116
rect 287 3096 289 3116
rect 301 3096 303 3116
rect 307 3096 311 3116
rect 315 3096 317 3116
rect 355 3096 357 3116
rect 361 3096 365 3116
rect 377 3096 379 3116
rect 383 3096 389 3116
rect 393 3096 395 3116
rect 407 3096 411 3116
rect 415 3096 421 3116
rect 425 3096 427 3116
rect 439 3096 441 3116
rect 255 3076 268 3096
rect 431 3076 441 3096
rect 445 3076 447 3116
rect 489 3076 491 3116
rect 495 3088 497 3116
rect 509 3088 511 3116
rect 495 3076 511 3088
rect 515 3076 517 3116
rect 529 3076 531 3116
rect 535 3076 537 3116
rect 591 3076 593 3116
rect 597 3076 603 3116
rect 607 3076 609 3116
rect 691 3076 693 3116
rect 697 3076 703 3116
rect 707 3076 709 3116
rect 763 3096 765 3116
rect 769 3096 771 3116
rect 783 3096 785 3116
rect 789 3096 791 3116
rect 831 3076 833 3116
rect 837 3076 843 3116
rect 847 3076 849 3116
rect 923 3076 925 3116
rect 929 3076 931 3116
rect 943 3076 945 3116
rect 949 3088 951 3116
rect 963 3088 965 3116
rect 949 3076 965 3088
rect 969 3076 971 3116
rect 1023 3076 1025 3116
rect 1029 3076 1031 3116
rect 1043 3076 1045 3116
rect 1049 3088 1051 3116
rect 1063 3088 1065 3116
rect 1049 3076 1065 3088
rect 1069 3076 1071 3116
rect 1123 3096 1125 3116
rect 1129 3096 1131 3116
rect 1143 3096 1145 3116
rect 1149 3096 1151 3116
rect 1203 3076 1205 3116
rect 1209 3076 1211 3116
rect 1223 3076 1225 3116
rect 1229 3088 1231 3116
rect 1243 3088 1245 3116
rect 1229 3076 1245 3088
rect 1249 3076 1251 3116
rect 1291 3076 1293 3116
rect 1297 3076 1303 3116
rect 1307 3076 1309 3116
rect 1383 3076 1385 3116
rect 1389 3076 1391 3116
rect 1431 3076 1433 3116
rect 1437 3076 1443 3116
rect 1447 3076 1449 3116
rect 1511 3076 1513 3116
rect 1517 3076 1523 3116
rect 1527 3076 1529 3116
rect 1589 3096 1591 3116
rect 1595 3096 1599 3116
rect 1611 3076 1613 3116
rect 1617 3076 1619 3116
rect 1669 3076 1671 3116
rect 1675 3088 1677 3116
rect 1689 3088 1691 3116
rect 1675 3076 1691 3088
rect 1695 3076 1697 3116
rect 1709 3076 1711 3116
rect 1715 3076 1717 3116
rect 1769 3076 1771 3116
rect 1775 3088 1777 3116
rect 1789 3088 1791 3116
rect 1775 3076 1791 3088
rect 1795 3076 1797 3116
rect 1809 3076 1811 3116
rect 1815 3076 1817 3116
rect 1869 3096 1871 3116
rect 1875 3096 1877 3116
rect 1889 3096 1891 3116
rect 1895 3096 1897 3116
rect 1952 3076 1954 3116
rect 1958 3076 1962 3116
rect 1966 3076 1968 3116
rect 1980 3096 1984 3116
rect 1988 3096 1990 3116
rect 2049 3096 2051 3116
rect 2055 3096 2057 3116
rect 2109 3076 2111 3116
rect 2115 3088 2117 3116
rect 2129 3088 2131 3116
rect 2115 3076 2131 3088
rect 2135 3076 2137 3116
rect 2149 3076 2151 3116
rect 2155 3076 2157 3116
rect 2209 3096 2211 3116
rect 2215 3096 2217 3116
rect 2229 3096 2231 3116
rect 2235 3096 2237 3116
rect 2311 3076 2313 3116
rect 2317 3076 2323 3116
rect 2327 3076 2329 3116
rect 2369 3076 2371 3116
rect 2375 3088 2377 3116
rect 2389 3088 2391 3116
rect 2375 3076 2391 3088
rect 2395 3076 2397 3116
rect 2409 3076 2411 3116
rect 2415 3076 2417 3116
rect 2469 3096 2471 3116
rect 2475 3096 2477 3116
rect 2529 3076 2531 3116
rect 2535 3088 2537 3116
rect 2549 3088 2551 3116
rect 2535 3076 2551 3088
rect 2555 3076 2557 3116
rect 2569 3076 2571 3116
rect 2575 3076 2577 3116
rect 2629 3096 2631 3116
rect 2635 3096 2639 3116
rect 2651 3076 2653 3116
rect 2657 3076 2659 3116
rect 2711 3076 2713 3116
rect 2717 3076 2723 3116
rect 2727 3076 2729 3116
rect 2793 3076 2795 3116
rect 2799 3096 2801 3116
rect 2813 3096 2815 3116
rect 2819 3096 2825 3116
rect 2829 3096 2833 3116
rect 2845 3096 2847 3116
rect 2851 3096 2857 3116
rect 2861 3096 2863 3116
rect 2875 3096 2879 3116
rect 2883 3096 2885 3116
rect 2923 3096 2925 3116
rect 2929 3096 2933 3116
rect 2937 3096 2939 3116
rect 2951 3096 2953 3116
rect 2957 3096 2963 3116
rect 2967 3096 2969 3116
rect 2981 3096 2985 3116
rect 2799 3076 2809 3096
rect 2972 3076 2985 3096
rect 2989 3076 2991 3116
rect 3043 3096 3045 3116
rect 3049 3096 3051 3116
rect 3063 3096 3065 3116
rect 3069 3096 3071 3116
rect 3130 3096 3132 3116
rect 3136 3096 3140 3116
rect 3152 3076 3154 3116
rect 3158 3076 3162 3116
rect 3166 3076 3168 3116
rect 3209 3096 3211 3116
rect 3215 3096 3217 3116
rect 3229 3096 3231 3116
rect 3235 3096 3237 3116
rect 3293 3076 3295 3116
rect 3299 3096 3301 3116
rect 3313 3096 3315 3116
rect 3319 3096 3325 3116
rect 3329 3096 3333 3116
rect 3345 3096 3347 3116
rect 3351 3096 3357 3116
rect 3361 3096 3363 3116
rect 3375 3096 3379 3116
rect 3383 3096 3385 3116
rect 3423 3096 3425 3116
rect 3429 3096 3433 3116
rect 3437 3096 3439 3116
rect 3451 3096 3453 3116
rect 3457 3096 3463 3116
rect 3467 3096 3469 3116
rect 3481 3096 3485 3116
rect 3299 3076 3309 3096
rect 3472 3076 3485 3096
rect 3489 3076 3491 3116
rect 3533 3076 3535 3116
rect 3539 3096 3541 3116
rect 3553 3096 3555 3116
rect 3559 3096 3565 3116
rect 3569 3096 3573 3116
rect 3585 3096 3587 3116
rect 3591 3096 3597 3116
rect 3601 3096 3603 3116
rect 3615 3096 3619 3116
rect 3623 3096 3625 3116
rect 3663 3096 3665 3116
rect 3669 3096 3673 3116
rect 3677 3096 3679 3116
rect 3691 3096 3693 3116
rect 3697 3096 3703 3116
rect 3707 3096 3709 3116
rect 3721 3096 3725 3116
rect 3539 3076 3549 3096
rect 3712 3076 3725 3096
rect 3729 3076 3731 3116
rect 3769 3096 3771 3116
rect 3775 3096 3777 3116
rect 3789 3096 3791 3116
rect 3795 3096 3797 3116
rect 3863 3076 3865 3116
rect 3869 3076 3871 3116
rect 3883 3076 3885 3116
rect 3889 3088 3891 3116
rect 3903 3088 3905 3116
rect 3889 3076 3905 3088
rect 3909 3076 3911 3116
rect 3963 3076 3965 3116
rect 3969 3076 3971 3116
rect 3983 3076 3985 3116
rect 3989 3088 3991 3116
rect 4003 3088 4005 3116
rect 3989 3076 4005 3088
rect 4009 3076 4011 3116
rect 4049 3076 4051 3116
rect 4055 3088 4057 3116
rect 4069 3088 4071 3116
rect 4055 3076 4071 3088
rect 4075 3076 4077 3116
rect 4089 3076 4091 3116
rect 4095 3076 4097 3116
rect 4149 3076 4151 3116
rect 4155 3088 4157 3116
rect 4169 3088 4171 3116
rect 4155 3076 4171 3088
rect 4175 3076 4177 3116
rect 4189 3076 4191 3116
rect 4195 3076 4197 3116
rect 4249 3096 4251 3116
rect 4255 3096 4257 3116
rect 4310 3056 4312 3116
rect 4316 3056 4320 3116
rect 4324 3056 4328 3116
rect 4332 3058 4334 3116
rect 4409 3076 4411 3116
rect 4415 3096 4419 3116
rect 4431 3096 4433 3116
rect 4437 3096 4443 3116
rect 4447 3096 4449 3116
rect 4461 3096 4463 3116
rect 4467 3096 4471 3116
rect 4475 3096 4477 3116
rect 4515 3096 4517 3116
rect 4521 3096 4525 3116
rect 4537 3096 4539 3116
rect 4543 3096 4549 3116
rect 4553 3096 4555 3116
rect 4567 3096 4571 3116
rect 4575 3096 4581 3116
rect 4585 3096 4587 3116
rect 4599 3096 4601 3116
rect 4415 3076 4428 3096
rect 4332 3056 4346 3058
rect 4591 3076 4601 3096
rect 4605 3076 4607 3116
rect 4649 3076 4651 3116
rect 4655 3088 4657 3116
rect 4669 3088 4671 3116
rect 4655 3076 4671 3088
rect 4675 3076 4677 3116
rect 4689 3076 4691 3116
rect 4695 3076 4697 3116
rect 43 2664 45 2684
rect 49 2664 51 2684
rect 103 2664 105 2704
rect 109 2664 111 2704
rect 123 2664 125 2704
rect 129 2692 145 2704
rect 129 2664 131 2692
rect 143 2664 145 2692
rect 149 2664 151 2704
rect 192 2664 194 2704
rect 198 2664 202 2704
rect 206 2664 208 2704
rect 220 2664 222 2704
rect 226 2664 230 2704
rect 234 2664 236 2704
rect 311 2664 313 2704
rect 317 2664 323 2704
rect 327 2664 329 2704
rect 389 2664 391 2704
rect 395 2664 401 2704
rect 405 2664 407 2704
rect 419 2664 421 2704
rect 425 2664 427 2704
rect 503 2664 505 2704
rect 509 2664 511 2704
rect 523 2664 525 2704
rect 529 2692 545 2704
rect 529 2664 531 2692
rect 543 2664 545 2692
rect 549 2664 551 2704
rect 591 2664 593 2704
rect 597 2664 603 2704
rect 607 2664 609 2704
rect 683 2664 685 2704
rect 689 2664 691 2704
rect 743 2664 745 2704
rect 749 2664 751 2704
rect 791 2664 793 2704
rect 797 2664 803 2704
rect 807 2664 809 2704
rect 869 2664 871 2704
rect 875 2664 881 2704
rect 885 2664 887 2704
rect 899 2664 901 2704
rect 905 2664 907 2704
rect 983 2664 985 2704
rect 989 2664 991 2704
rect 1003 2664 1005 2704
rect 1009 2692 1025 2704
rect 1009 2664 1011 2692
rect 1023 2664 1025 2692
rect 1029 2664 1031 2704
rect 1071 2664 1073 2704
rect 1077 2664 1083 2704
rect 1087 2664 1089 2704
rect 1163 2664 1165 2704
rect 1169 2664 1171 2704
rect 1183 2664 1185 2704
rect 1189 2692 1205 2704
rect 1189 2664 1191 2692
rect 1203 2664 1205 2692
rect 1209 2664 1211 2704
rect 1249 2664 1251 2704
rect 1255 2684 1268 2704
rect 1431 2684 1441 2704
rect 1255 2664 1259 2684
rect 1271 2664 1273 2684
rect 1277 2664 1283 2684
rect 1287 2664 1289 2684
rect 1301 2664 1303 2684
rect 1307 2664 1311 2684
rect 1315 2664 1317 2684
rect 1355 2664 1357 2684
rect 1361 2664 1365 2684
rect 1377 2664 1379 2684
rect 1383 2664 1389 2684
rect 1393 2664 1395 2684
rect 1407 2664 1411 2684
rect 1415 2664 1421 2684
rect 1425 2664 1427 2684
rect 1439 2664 1441 2684
rect 1445 2664 1447 2704
rect 1501 2664 1503 2704
rect 1507 2664 1509 2704
rect 1521 2664 1525 2684
rect 1529 2664 1531 2684
rect 1573 2664 1575 2704
rect 1579 2684 1589 2704
rect 1752 2684 1765 2704
rect 1579 2664 1581 2684
rect 1593 2664 1595 2684
rect 1599 2664 1605 2684
rect 1609 2664 1613 2684
rect 1625 2664 1627 2684
rect 1631 2664 1637 2684
rect 1641 2664 1643 2684
rect 1655 2664 1659 2684
rect 1663 2664 1665 2684
rect 1703 2664 1705 2684
rect 1709 2664 1713 2684
rect 1717 2664 1719 2684
rect 1731 2664 1733 2684
rect 1737 2664 1743 2684
rect 1747 2664 1749 2684
rect 1761 2664 1765 2684
rect 1769 2664 1771 2704
rect 1809 2664 1811 2704
rect 1815 2692 1831 2704
rect 1815 2664 1817 2692
rect 1829 2664 1831 2692
rect 1835 2664 1837 2704
rect 1849 2664 1851 2704
rect 1855 2664 1857 2704
rect 1909 2664 1911 2684
rect 1915 2664 1917 2684
rect 1969 2664 1971 2704
rect 1975 2694 1991 2704
rect 1975 2664 1977 2694
rect 1989 2664 1991 2694
rect 1995 2664 1997 2704
rect 2009 2664 2011 2704
rect 2015 2676 2017 2704
rect 2029 2676 2031 2704
rect 2015 2664 2031 2676
rect 2035 2664 2037 2704
rect 2103 2664 2105 2684
rect 2109 2664 2111 2684
rect 2123 2664 2125 2684
rect 2129 2664 2131 2684
rect 2183 2664 2185 2684
rect 2189 2664 2191 2684
rect 2203 2664 2205 2684
rect 2209 2664 2211 2684
rect 2263 2664 2265 2684
rect 2269 2664 2271 2684
rect 2283 2664 2285 2684
rect 2289 2664 2291 2684
rect 2329 2664 2331 2684
rect 2335 2664 2337 2684
rect 2403 2664 2405 2684
rect 2409 2664 2411 2684
rect 2423 2664 2425 2684
rect 2429 2664 2431 2684
rect 2469 2664 2471 2684
rect 2475 2664 2477 2684
rect 2529 2664 2531 2704
rect 2535 2664 2541 2704
rect 2545 2664 2547 2704
rect 2559 2664 2561 2704
rect 2565 2664 2567 2704
rect 2629 2664 2631 2704
rect 2635 2692 2651 2704
rect 2635 2664 2637 2692
rect 2649 2664 2651 2692
rect 2655 2664 2657 2704
rect 2669 2664 2671 2704
rect 2675 2664 2677 2704
rect 2729 2664 2731 2704
rect 2735 2692 2751 2704
rect 2735 2664 2737 2692
rect 2749 2664 2751 2692
rect 2755 2664 2757 2704
rect 2769 2664 2771 2704
rect 2775 2664 2777 2704
rect 2831 2664 2833 2704
rect 2837 2664 2843 2704
rect 2847 2664 2849 2704
rect 2913 2664 2915 2704
rect 2919 2684 2929 2704
rect 3092 2684 3105 2704
rect 2919 2664 2921 2684
rect 2933 2664 2935 2684
rect 2939 2664 2945 2684
rect 2949 2664 2953 2684
rect 2965 2664 2967 2684
rect 2971 2664 2977 2684
rect 2981 2664 2983 2684
rect 2995 2664 2999 2684
rect 3003 2664 3005 2684
rect 3043 2664 3045 2684
rect 3049 2664 3053 2684
rect 3057 2664 3059 2684
rect 3071 2664 3073 2684
rect 3077 2664 3083 2684
rect 3087 2664 3089 2684
rect 3101 2664 3105 2684
rect 3109 2664 3111 2704
rect 3153 2664 3155 2704
rect 3159 2684 3169 2704
rect 3332 2684 3345 2704
rect 3159 2664 3161 2684
rect 3173 2664 3175 2684
rect 3179 2664 3185 2684
rect 3189 2664 3193 2684
rect 3205 2664 3207 2684
rect 3211 2664 3217 2684
rect 3221 2664 3223 2684
rect 3235 2664 3239 2684
rect 3243 2664 3245 2684
rect 3283 2664 3285 2684
rect 3289 2664 3293 2684
rect 3297 2664 3299 2684
rect 3311 2664 3313 2684
rect 3317 2664 3323 2684
rect 3327 2664 3329 2684
rect 3341 2664 3345 2684
rect 3349 2664 3351 2704
rect 3403 2664 3405 2684
rect 3409 2664 3411 2684
rect 3463 2664 3465 2684
rect 3469 2664 3471 2684
rect 3483 2664 3485 2684
rect 3489 2664 3491 2684
rect 3543 2664 3545 2704
rect 3549 2664 3551 2704
rect 3593 2664 3595 2704
rect 3599 2684 3609 2704
rect 3772 2684 3785 2704
rect 3599 2664 3601 2684
rect 3613 2664 3615 2684
rect 3619 2664 3625 2684
rect 3629 2664 3633 2684
rect 3645 2664 3647 2684
rect 3651 2664 3657 2684
rect 3661 2664 3663 2684
rect 3675 2664 3679 2684
rect 3683 2664 3685 2684
rect 3723 2664 3725 2684
rect 3729 2664 3733 2684
rect 3737 2664 3739 2684
rect 3751 2664 3753 2684
rect 3757 2664 3763 2684
rect 3767 2664 3769 2684
rect 3781 2664 3785 2684
rect 3789 2664 3791 2704
rect 3864 2664 3866 2704
rect 3870 2664 3874 2704
rect 3878 2664 3880 2704
rect 3892 2664 3894 2704
rect 3898 2664 3902 2704
rect 3906 2664 3908 2704
rect 3963 2664 3965 2684
rect 3969 2664 3971 2684
rect 3983 2664 3985 2684
rect 3989 2664 3991 2684
rect 4029 2664 4031 2704
rect 4035 2692 4051 2704
rect 4035 2664 4037 2692
rect 4049 2664 4051 2692
rect 4055 2664 4057 2704
rect 4069 2664 4071 2704
rect 4075 2664 4077 2704
rect 4143 2664 4145 2704
rect 4149 2664 4151 2704
rect 4163 2664 4165 2704
rect 4169 2692 4185 2704
rect 4169 2664 4171 2692
rect 4183 2664 4185 2692
rect 4189 2664 4191 2704
rect 4229 2664 4231 2684
rect 4235 2664 4237 2684
rect 4249 2664 4251 2684
rect 4255 2664 4257 2684
rect 4313 2664 4315 2704
rect 4319 2684 4329 2704
rect 4492 2684 4505 2704
rect 4319 2664 4321 2684
rect 4333 2664 4335 2684
rect 4339 2664 4345 2684
rect 4349 2664 4353 2684
rect 4365 2664 4367 2684
rect 4371 2664 4377 2684
rect 4381 2664 4383 2684
rect 4395 2664 4399 2684
rect 4403 2664 4405 2684
rect 4443 2664 4445 2684
rect 4449 2664 4453 2684
rect 4457 2664 4459 2684
rect 4471 2664 4473 2684
rect 4477 2664 4483 2684
rect 4487 2664 4489 2684
rect 4501 2664 4505 2684
rect 4509 2664 4511 2704
rect 4549 2664 4551 2704
rect 4555 2692 4571 2704
rect 4555 2664 4557 2692
rect 4569 2664 4571 2692
rect 4575 2664 4577 2704
rect 4589 2664 4591 2704
rect 4595 2664 4597 2704
rect 4651 2664 4653 2704
rect 4657 2664 4663 2704
rect 4667 2664 4669 2704
rect 30 2576 32 2636
rect 36 2576 40 2636
rect 44 2576 48 2636
rect 52 2578 54 2636
rect 132 2596 134 2636
rect 138 2596 142 2636
rect 146 2596 148 2636
rect 160 2616 164 2636
rect 168 2616 170 2636
rect 243 2616 245 2636
rect 249 2616 251 2636
rect 52 2576 66 2578
rect 313 2596 315 2636
rect 319 2596 321 2636
rect 333 2596 335 2636
rect 339 2596 345 2636
rect 349 2596 351 2636
rect 410 2616 412 2636
rect 416 2616 420 2636
rect 432 2596 434 2636
rect 438 2596 442 2636
rect 446 2596 448 2636
rect 526 2578 528 2636
rect 514 2576 528 2578
rect 532 2576 536 2636
rect 540 2576 544 2636
rect 548 2576 550 2636
rect 603 2596 605 2636
rect 609 2596 611 2636
rect 623 2596 625 2636
rect 629 2608 631 2636
rect 643 2608 645 2636
rect 629 2596 645 2608
rect 649 2596 651 2636
rect 703 2596 705 2636
rect 709 2596 711 2636
rect 771 2596 773 2636
rect 777 2596 783 2636
rect 787 2596 789 2636
rect 866 2578 868 2636
rect 854 2576 868 2578
rect 872 2576 876 2636
rect 880 2576 884 2636
rect 888 2576 890 2636
rect 943 2596 945 2636
rect 949 2596 951 2636
rect 963 2596 965 2636
rect 969 2608 971 2636
rect 983 2608 985 2636
rect 969 2596 985 2608
rect 989 2596 991 2636
rect 1031 2596 1033 2636
rect 1037 2596 1043 2636
rect 1047 2596 1049 2636
rect 1146 2578 1148 2636
rect 1134 2576 1148 2578
rect 1152 2576 1156 2636
rect 1160 2576 1164 2636
rect 1168 2576 1170 2636
rect 1223 2616 1225 2636
rect 1229 2616 1231 2636
rect 1283 2596 1285 2636
rect 1289 2596 1291 2636
rect 1303 2596 1305 2636
rect 1309 2608 1311 2636
rect 1323 2608 1325 2636
rect 1309 2596 1325 2608
rect 1329 2596 1331 2636
rect 1371 2596 1373 2636
rect 1377 2596 1383 2636
rect 1387 2596 1389 2636
rect 1449 2596 1451 2636
rect 1455 2596 1457 2636
rect 1531 2596 1533 2636
rect 1537 2596 1543 2636
rect 1547 2596 1549 2636
rect 1593 2596 1595 2636
rect 1599 2616 1601 2636
rect 1613 2616 1615 2636
rect 1619 2616 1625 2636
rect 1629 2616 1633 2636
rect 1645 2616 1647 2636
rect 1651 2616 1657 2636
rect 1661 2616 1663 2636
rect 1675 2616 1679 2636
rect 1683 2616 1685 2636
rect 1723 2616 1725 2636
rect 1729 2616 1733 2636
rect 1737 2616 1739 2636
rect 1751 2616 1753 2636
rect 1757 2616 1763 2636
rect 1767 2616 1769 2636
rect 1781 2616 1785 2636
rect 1599 2596 1609 2616
rect 1772 2596 1785 2616
rect 1789 2596 1791 2636
rect 1831 2596 1833 2636
rect 1837 2596 1843 2636
rect 1847 2596 1849 2636
rect 1911 2596 1913 2636
rect 1917 2596 1923 2636
rect 1927 2596 1929 2636
rect 1990 2576 1992 2636
rect 1996 2576 2000 2636
rect 2004 2576 2008 2636
rect 2012 2578 2014 2636
rect 2089 2616 2091 2636
rect 2095 2616 2097 2636
rect 2109 2616 2111 2636
rect 2115 2616 2117 2636
rect 2183 2616 2185 2636
rect 2189 2616 2191 2636
rect 2243 2616 2245 2636
rect 2249 2616 2251 2636
rect 2263 2616 2265 2636
rect 2269 2616 2271 2636
rect 2323 2616 2325 2636
rect 2329 2616 2331 2636
rect 2012 2576 2026 2578
rect 2383 2596 2385 2636
rect 2389 2596 2391 2636
rect 2403 2596 2405 2636
rect 2409 2608 2411 2636
rect 2423 2608 2425 2636
rect 2409 2596 2425 2608
rect 2429 2596 2431 2636
rect 2469 2616 2471 2636
rect 2475 2616 2477 2636
rect 2489 2616 2491 2636
rect 2495 2616 2497 2636
rect 2549 2596 2551 2636
rect 2555 2596 2561 2636
rect 2565 2596 2567 2636
rect 2579 2596 2581 2636
rect 2585 2596 2587 2636
rect 2649 2596 2651 2636
rect 2655 2608 2657 2636
rect 2669 2608 2671 2636
rect 2655 2596 2671 2608
rect 2675 2596 2677 2636
rect 2689 2596 2691 2636
rect 2695 2596 2697 2636
rect 2771 2596 2773 2636
rect 2777 2596 2783 2636
rect 2787 2596 2789 2636
rect 2829 2616 2831 2636
rect 2835 2616 2837 2636
rect 2849 2616 2851 2636
rect 2855 2616 2857 2636
rect 2869 2616 2871 2636
rect 2859 2596 2871 2616
rect 2875 2596 2877 2636
rect 2931 2596 2933 2636
rect 2937 2596 2943 2636
rect 2947 2596 2949 2636
rect 3009 2616 3011 2636
rect 3015 2616 3019 2636
rect 3031 2596 3033 2636
rect 3037 2596 3039 2636
rect 3089 2596 3091 2636
rect 3095 2608 3097 2636
rect 3109 2608 3111 2636
rect 3095 2596 3111 2608
rect 3115 2596 3117 2636
rect 3129 2596 3131 2636
rect 3135 2596 3137 2636
rect 3201 2596 3203 2636
rect 3207 2596 3209 2636
rect 3221 2616 3225 2636
rect 3229 2616 3231 2636
rect 3291 2596 3293 2636
rect 3297 2596 3303 2636
rect 3307 2596 3309 2636
rect 3352 2596 3354 2636
rect 3358 2596 3362 2636
rect 3366 2596 3368 2636
rect 3380 2596 3382 2636
rect 3386 2596 3390 2636
rect 3394 2596 3396 2636
rect 3469 2616 3471 2636
rect 3475 2616 3479 2636
rect 3491 2596 3493 2636
rect 3497 2596 3499 2636
rect 3561 2596 3563 2636
rect 3567 2596 3569 2636
rect 3581 2616 3585 2636
rect 3589 2616 3591 2636
rect 3633 2596 3635 2636
rect 3639 2616 3641 2636
rect 3653 2616 3655 2636
rect 3659 2616 3665 2636
rect 3669 2616 3673 2636
rect 3685 2616 3687 2636
rect 3691 2616 3697 2636
rect 3701 2616 3703 2636
rect 3715 2616 3719 2636
rect 3723 2616 3725 2636
rect 3763 2616 3765 2636
rect 3769 2616 3773 2636
rect 3777 2616 3779 2636
rect 3791 2616 3793 2636
rect 3797 2616 3803 2636
rect 3807 2616 3809 2636
rect 3821 2616 3825 2636
rect 3639 2596 3649 2616
rect 3812 2596 3825 2616
rect 3829 2596 3831 2636
rect 3890 2616 3892 2636
rect 3896 2616 3900 2636
rect 3912 2596 3914 2636
rect 3918 2596 3922 2636
rect 3926 2596 3928 2636
rect 3969 2616 3971 2636
rect 3975 2616 3977 2636
rect 3989 2616 3991 2636
rect 3995 2616 3997 2636
rect 4049 2596 4051 2636
rect 4055 2596 4057 2636
rect 4069 2596 4071 2636
rect 4075 2596 4077 2636
rect 4089 2596 4091 2636
rect 4095 2596 4097 2636
rect 4109 2596 4111 2636
rect 4115 2596 4117 2636
rect 4129 2596 4131 2636
rect 4135 2596 4137 2636
rect 4149 2596 4151 2636
rect 4155 2596 4157 2636
rect 4169 2596 4171 2636
rect 4175 2596 4177 2636
rect 4189 2596 4191 2636
rect 4195 2596 4197 2636
rect 4253 2596 4255 2636
rect 4259 2616 4261 2636
rect 4273 2616 4275 2636
rect 4279 2616 4285 2636
rect 4289 2616 4293 2636
rect 4305 2616 4307 2636
rect 4311 2616 4317 2636
rect 4321 2616 4323 2636
rect 4335 2616 4339 2636
rect 4343 2616 4345 2636
rect 4383 2616 4385 2636
rect 4389 2616 4393 2636
rect 4397 2616 4399 2636
rect 4411 2616 4413 2636
rect 4417 2616 4423 2636
rect 4427 2616 4429 2636
rect 4441 2616 4445 2636
rect 4259 2596 4269 2616
rect 4432 2596 4445 2616
rect 4449 2596 4451 2636
rect 4489 2596 4491 2636
rect 4495 2608 4497 2636
rect 4509 2608 4511 2636
rect 4495 2596 4511 2608
rect 4515 2596 4517 2636
rect 4529 2596 4531 2636
rect 4535 2596 4537 2636
rect 4591 2596 4593 2636
rect 4597 2596 4603 2636
rect 4607 2596 4609 2636
rect 4671 2596 4673 2636
rect 4677 2596 4683 2636
rect 4687 2596 4689 2636
rect 54 2242 68 2244
rect 66 2184 68 2242
rect 72 2184 76 2244
rect 80 2184 84 2244
rect 88 2184 90 2244
rect 143 2184 145 2224
rect 149 2184 151 2224
rect 163 2184 165 2224
rect 169 2212 185 2224
rect 169 2184 171 2212
rect 183 2184 185 2212
rect 189 2184 191 2224
rect 229 2184 231 2224
rect 235 2212 251 2224
rect 235 2184 237 2212
rect 249 2184 251 2212
rect 255 2184 257 2224
rect 269 2184 271 2224
rect 275 2184 277 2224
rect 330 2184 332 2244
rect 336 2184 340 2244
rect 344 2184 348 2244
rect 352 2242 366 2244
rect 352 2184 354 2242
rect 432 2184 434 2224
rect 438 2184 442 2224
rect 446 2184 448 2224
rect 460 2184 464 2204
rect 468 2184 470 2204
rect 529 2184 531 2224
rect 535 2212 551 2224
rect 535 2184 537 2212
rect 549 2184 551 2212
rect 555 2184 557 2224
rect 569 2184 571 2224
rect 575 2184 577 2224
rect 650 2184 652 2204
rect 656 2184 660 2204
rect 672 2184 674 2224
rect 678 2184 682 2224
rect 686 2184 688 2224
rect 729 2184 731 2204
rect 735 2184 737 2204
rect 813 2184 815 2224
rect 819 2184 821 2224
rect 833 2184 835 2224
rect 839 2184 845 2224
rect 849 2184 851 2224
rect 891 2184 893 2224
rect 897 2184 903 2224
rect 907 2184 909 2224
rect 969 2184 971 2224
rect 975 2184 981 2224
rect 985 2184 987 2224
rect 999 2184 1001 2224
rect 1005 2184 1007 2224
rect 1083 2184 1085 2224
rect 1089 2184 1091 2224
rect 1103 2184 1105 2224
rect 1109 2212 1125 2224
rect 1109 2184 1111 2212
rect 1123 2184 1125 2212
rect 1129 2184 1131 2224
rect 1183 2184 1185 2224
rect 1189 2184 1191 2224
rect 1203 2184 1205 2224
rect 1209 2212 1225 2224
rect 1209 2184 1211 2212
rect 1223 2184 1225 2212
rect 1229 2184 1231 2224
rect 1273 2184 1275 2224
rect 1279 2204 1289 2224
rect 1452 2204 1465 2224
rect 1279 2184 1281 2204
rect 1293 2184 1295 2204
rect 1299 2184 1305 2204
rect 1309 2184 1313 2204
rect 1325 2184 1327 2204
rect 1331 2184 1337 2204
rect 1341 2184 1343 2204
rect 1355 2184 1359 2204
rect 1363 2184 1365 2204
rect 1403 2184 1405 2204
rect 1409 2184 1413 2204
rect 1417 2184 1419 2204
rect 1431 2184 1433 2204
rect 1437 2184 1443 2204
rect 1447 2184 1449 2204
rect 1461 2184 1465 2204
rect 1469 2184 1471 2224
rect 1523 2184 1525 2224
rect 1529 2184 1531 2224
rect 1543 2184 1545 2224
rect 1549 2212 1565 2224
rect 1549 2184 1551 2212
rect 1563 2184 1565 2212
rect 1569 2184 1571 2224
rect 1613 2184 1615 2224
rect 1619 2204 1629 2224
rect 1792 2204 1805 2224
rect 1619 2184 1621 2204
rect 1633 2184 1635 2204
rect 1639 2184 1645 2204
rect 1649 2184 1653 2204
rect 1665 2184 1667 2204
rect 1671 2184 1677 2204
rect 1681 2184 1683 2204
rect 1695 2184 1699 2204
rect 1703 2184 1705 2204
rect 1743 2184 1745 2204
rect 1749 2184 1753 2204
rect 1757 2184 1759 2204
rect 1771 2184 1773 2204
rect 1777 2184 1783 2204
rect 1787 2184 1789 2204
rect 1801 2184 1805 2204
rect 1809 2184 1811 2224
rect 1863 2184 1865 2204
rect 1869 2184 1871 2204
rect 1923 2184 1925 2204
rect 1929 2184 1931 2204
rect 1969 2184 1971 2224
rect 1975 2212 1991 2224
rect 1975 2184 1977 2212
rect 1989 2184 1991 2212
rect 1995 2184 1997 2224
rect 2009 2184 2011 2224
rect 2015 2184 2017 2224
rect 2073 2184 2075 2224
rect 2079 2204 2089 2224
rect 2252 2204 2265 2224
rect 2079 2184 2081 2204
rect 2093 2184 2095 2204
rect 2099 2184 2105 2204
rect 2109 2184 2113 2204
rect 2125 2184 2127 2204
rect 2131 2184 2137 2204
rect 2141 2184 2143 2204
rect 2155 2184 2159 2204
rect 2163 2184 2165 2204
rect 2203 2184 2205 2204
rect 2209 2184 2213 2204
rect 2217 2184 2219 2204
rect 2231 2184 2233 2204
rect 2237 2184 2243 2204
rect 2247 2184 2249 2204
rect 2261 2184 2265 2204
rect 2269 2184 2271 2224
rect 2330 2184 2332 2204
rect 2336 2184 2340 2204
rect 2352 2184 2354 2224
rect 2358 2184 2362 2224
rect 2366 2184 2368 2224
rect 2430 2184 2432 2204
rect 2436 2184 2440 2204
rect 2452 2184 2454 2224
rect 2458 2184 2462 2224
rect 2466 2184 2468 2224
rect 2510 2184 2512 2244
rect 2516 2184 2520 2244
rect 2524 2184 2528 2244
rect 2532 2242 2546 2244
rect 2532 2184 2534 2242
rect 2609 2184 2611 2224
rect 2615 2184 2621 2224
rect 2625 2184 2627 2224
rect 2639 2184 2641 2224
rect 2645 2184 2647 2224
rect 2709 2184 2711 2224
rect 2715 2204 2728 2224
rect 2891 2204 2901 2224
rect 2715 2184 2719 2204
rect 2731 2184 2733 2204
rect 2737 2184 2743 2204
rect 2747 2184 2749 2204
rect 2761 2184 2763 2204
rect 2767 2184 2771 2204
rect 2775 2184 2777 2204
rect 2815 2184 2817 2204
rect 2821 2184 2825 2204
rect 2837 2184 2839 2204
rect 2843 2184 2849 2204
rect 2853 2184 2855 2204
rect 2867 2184 2871 2204
rect 2875 2184 2881 2204
rect 2885 2184 2887 2204
rect 2899 2184 2901 2204
rect 2905 2184 2907 2224
rect 2963 2184 2965 2224
rect 2969 2184 2971 2224
rect 2983 2184 2985 2224
rect 2989 2212 3005 2224
rect 2989 2184 2991 2212
rect 3003 2184 3005 2212
rect 3009 2184 3011 2224
rect 3063 2184 3065 2224
rect 3069 2184 3071 2224
rect 3083 2184 3085 2224
rect 3089 2212 3105 2224
rect 3089 2184 3091 2212
rect 3103 2184 3105 2212
rect 3109 2184 3111 2224
rect 3149 2184 3151 2224
rect 3155 2212 3171 2224
rect 3155 2184 3157 2212
rect 3169 2184 3171 2212
rect 3175 2184 3177 2224
rect 3189 2184 3191 2224
rect 3195 2184 3197 2224
rect 3249 2184 3251 2224
rect 3255 2204 3268 2224
rect 3431 2204 3441 2224
rect 3255 2184 3259 2204
rect 3271 2184 3273 2204
rect 3277 2184 3283 2204
rect 3287 2184 3289 2204
rect 3301 2184 3303 2204
rect 3307 2184 3311 2204
rect 3315 2184 3317 2204
rect 3355 2184 3357 2204
rect 3361 2184 3365 2204
rect 3377 2184 3379 2204
rect 3383 2184 3389 2204
rect 3393 2184 3395 2204
rect 3407 2184 3411 2204
rect 3415 2184 3421 2204
rect 3425 2184 3427 2204
rect 3439 2184 3441 2204
rect 3445 2184 3447 2224
rect 3503 2184 3505 2224
rect 3509 2184 3511 2224
rect 3523 2184 3525 2224
rect 3529 2212 3545 2224
rect 3529 2184 3531 2212
rect 3543 2184 3545 2212
rect 3549 2184 3551 2224
rect 3699 2204 3711 2224
rect 3603 2184 3605 2204
rect 3609 2184 3611 2204
rect 3623 2184 3625 2204
rect 3629 2184 3631 2204
rect 3669 2184 3671 2204
rect 3675 2184 3677 2204
rect 3689 2184 3691 2204
rect 3695 2184 3697 2204
rect 3709 2184 3711 2204
rect 3715 2184 3717 2224
rect 3791 2184 3793 2224
rect 3797 2184 3803 2224
rect 3807 2184 3809 2224
rect 3884 2184 3886 2224
rect 3890 2184 3894 2224
rect 3898 2184 3900 2224
rect 3912 2184 3914 2224
rect 3918 2184 3922 2224
rect 3926 2184 3928 2224
rect 4004 2184 4006 2224
rect 4010 2184 4014 2224
rect 4018 2184 4020 2224
rect 4032 2184 4034 2224
rect 4038 2184 4042 2224
rect 4046 2184 4048 2224
rect 4093 2184 4095 2224
rect 4099 2204 4109 2224
rect 4272 2204 4285 2224
rect 4099 2184 4101 2204
rect 4113 2184 4115 2204
rect 4119 2184 4125 2204
rect 4129 2184 4133 2204
rect 4145 2184 4147 2204
rect 4151 2184 4157 2204
rect 4161 2184 4163 2204
rect 4175 2184 4179 2204
rect 4183 2184 4185 2204
rect 4223 2184 4225 2204
rect 4229 2184 4233 2204
rect 4237 2184 4239 2204
rect 4251 2184 4253 2204
rect 4257 2184 4263 2204
rect 4267 2184 4269 2204
rect 4281 2184 4285 2204
rect 4289 2184 4291 2224
rect 4329 2184 4331 2224
rect 4335 2204 4348 2224
rect 4511 2204 4521 2224
rect 4335 2184 4339 2204
rect 4351 2184 4353 2204
rect 4357 2184 4363 2204
rect 4367 2184 4369 2204
rect 4381 2184 4383 2204
rect 4387 2184 4391 2204
rect 4395 2184 4397 2204
rect 4435 2184 4437 2204
rect 4441 2184 4445 2204
rect 4457 2184 4459 2204
rect 4463 2184 4469 2204
rect 4473 2184 4475 2204
rect 4487 2184 4491 2204
rect 4495 2184 4501 2204
rect 4505 2184 4507 2204
rect 4519 2184 4521 2204
rect 4525 2184 4527 2224
rect 4569 2184 4571 2224
rect 4575 2212 4591 2224
rect 4575 2184 4577 2212
rect 4589 2184 4591 2212
rect 4595 2184 4597 2224
rect 4609 2184 4611 2224
rect 4615 2184 4617 2224
rect 4671 2184 4673 2224
rect 4677 2184 4683 2224
rect 4687 2184 4689 2224
rect 41 2116 43 2156
rect 47 2116 49 2156
rect 61 2136 65 2156
rect 69 2136 71 2156
rect 123 2116 125 2156
rect 129 2116 131 2156
rect 143 2116 145 2156
rect 149 2128 151 2156
rect 163 2128 165 2156
rect 149 2116 165 2128
rect 169 2116 171 2156
rect 246 2098 248 2156
rect 234 2096 248 2098
rect 252 2096 256 2156
rect 260 2096 264 2156
rect 268 2096 270 2156
rect 312 2116 314 2156
rect 318 2116 322 2156
rect 326 2116 328 2156
rect 340 2136 344 2156
rect 348 2136 350 2156
rect 412 2116 414 2156
rect 418 2116 422 2156
rect 426 2116 428 2156
rect 440 2136 444 2156
rect 448 2136 450 2156
rect 510 2096 512 2156
rect 516 2096 520 2156
rect 524 2096 528 2156
rect 532 2098 534 2156
rect 532 2096 546 2098
rect 610 2096 612 2156
rect 616 2096 620 2156
rect 624 2096 628 2156
rect 632 2098 634 2156
rect 712 2116 714 2156
rect 718 2116 722 2156
rect 726 2116 728 2156
rect 740 2136 744 2156
rect 748 2136 750 2156
rect 632 2096 646 2098
rect 823 2116 825 2156
rect 829 2116 831 2156
rect 843 2116 845 2156
rect 849 2128 851 2156
rect 863 2128 865 2156
rect 849 2116 865 2128
rect 869 2116 871 2156
rect 910 2096 912 2156
rect 916 2096 920 2156
rect 924 2096 928 2156
rect 932 2098 934 2156
rect 932 2096 946 2098
rect 1010 2096 1012 2156
rect 1016 2096 1020 2156
rect 1024 2096 1028 2156
rect 1032 2098 1034 2156
rect 1032 2096 1046 2098
rect 1110 2096 1112 2156
rect 1116 2096 1120 2156
rect 1124 2096 1128 2156
rect 1132 2098 1134 2156
rect 1212 2116 1214 2156
rect 1218 2116 1222 2156
rect 1226 2116 1228 2156
rect 1240 2136 1244 2156
rect 1248 2136 1250 2156
rect 1309 2136 1311 2156
rect 1315 2136 1317 2156
rect 1329 2136 1331 2156
rect 1335 2136 1337 2156
rect 1132 2096 1146 2098
rect 1411 2116 1413 2156
rect 1417 2116 1423 2156
rect 1427 2116 1429 2156
rect 1491 2116 1493 2156
rect 1497 2116 1503 2156
rect 1507 2116 1509 2156
rect 1551 2116 1553 2156
rect 1557 2116 1563 2156
rect 1567 2116 1569 2156
rect 1643 2116 1645 2156
rect 1649 2116 1651 2156
rect 1663 2116 1665 2156
rect 1669 2128 1671 2156
rect 1683 2128 1685 2156
rect 1669 2116 1685 2128
rect 1689 2116 1691 2156
rect 1732 2116 1734 2156
rect 1738 2116 1742 2156
rect 1746 2116 1748 2156
rect 1760 2136 1764 2156
rect 1768 2136 1770 2156
rect 1829 2136 1831 2156
rect 1835 2136 1837 2156
rect 1849 2136 1851 2156
rect 1855 2136 1857 2156
rect 1923 2116 1925 2156
rect 1929 2116 1931 2156
rect 1943 2116 1945 2156
rect 1949 2128 1951 2156
rect 1963 2128 1965 2156
rect 1949 2116 1965 2128
rect 1969 2116 1971 2156
rect 2009 2116 2011 2156
rect 2015 2128 2017 2156
rect 2029 2128 2031 2156
rect 2015 2116 2031 2128
rect 2035 2116 2037 2156
rect 2049 2116 2051 2156
rect 2055 2116 2057 2156
rect 2123 2116 2125 2156
rect 2129 2116 2131 2156
rect 2143 2116 2145 2156
rect 2149 2128 2151 2156
rect 2163 2128 2165 2156
rect 2149 2116 2165 2128
rect 2169 2116 2171 2156
rect 2223 2116 2225 2156
rect 2229 2116 2231 2156
rect 2243 2116 2245 2156
rect 2249 2116 2251 2156
rect 2263 2116 2265 2156
rect 2269 2116 2271 2156
rect 2283 2116 2285 2156
rect 2289 2116 2291 2156
rect 2303 2116 2305 2156
rect 2309 2116 2311 2156
rect 2323 2116 2325 2156
rect 2329 2116 2331 2156
rect 2343 2116 2345 2156
rect 2349 2116 2351 2156
rect 2363 2116 2365 2156
rect 2369 2116 2371 2156
rect 2411 2116 2413 2156
rect 2417 2116 2423 2156
rect 2427 2116 2429 2156
rect 2513 2116 2515 2156
rect 2519 2116 2521 2156
rect 2533 2116 2535 2156
rect 2539 2116 2545 2156
rect 2549 2116 2551 2156
rect 2589 2136 2591 2156
rect 2595 2136 2597 2156
rect 2609 2136 2611 2156
rect 2615 2136 2617 2156
rect 2629 2136 2631 2156
rect 2619 2116 2631 2136
rect 2635 2116 2637 2156
rect 2711 2116 2713 2156
rect 2717 2116 2723 2156
rect 2727 2116 2729 2156
rect 2771 2116 2773 2156
rect 2777 2116 2783 2156
rect 2787 2116 2789 2156
rect 2853 2116 2855 2156
rect 2859 2136 2861 2156
rect 2873 2136 2875 2156
rect 2879 2136 2885 2156
rect 2889 2136 2893 2156
rect 2905 2136 2907 2156
rect 2911 2136 2917 2156
rect 2921 2136 2923 2156
rect 2935 2136 2939 2156
rect 2943 2136 2945 2156
rect 2983 2136 2985 2156
rect 2989 2136 2993 2156
rect 2997 2136 2999 2156
rect 3011 2136 3013 2156
rect 3017 2136 3023 2156
rect 3027 2136 3029 2156
rect 3041 2136 3045 2156
rect 2859 2116 2869 2136
rect 3032 2116 3045 2136
rect 3049 2116 3051 2156
rect 3110 2136 3112 2156
rect 3116 2136 3120 2156
rect 3132 2116 3134 2156
rect 3138 2116 3142 2156
rect 3146 2116 3148 2156
rect 3189 2136 3191 2156
rect 3195 2136 3197 2156
rect 3209 2136 3211 2156
rect 3215 2136 3217 2156
rect 3304 2116 3306 2156
rect 3310 2116 3314 2156
rect 3318 2116 3320 2156
rect 3332 2116 3334 2156
rect 3338 2116 3342 2156
rect 3346 2116 3348 2156
rect 3393 2116 3395 2156
rect 3399 2136 3401 2156
rect 3413 2136 3415 2156
rect 3419 2136 3425 2156
rect 3429 2136 3433 2156
rect 3445 2136 3447 2156
rect 3451 2136 3457 2156
rect 3461 2136 3463 2156
rect 3475 2136 3479 2156
rect 3483 2136 3485 2156
rect 3523 2136 3525 2156
rect 3529 2136 3533 2156
rect 3537 2136 3539 2156
rect 3551 2136 3553 2156
rect 3557 2136 3563 2156
rect 3567 2136 3569 2156
rect 3581 2136 3585 2156
rect 3399 2116 3409 2136
rect 3572 2116 3585 2136
rect 3589 2116 3591 2156
rect 3629 2116 3631 2156
rect 3635 2128 3637 2156
rect 3649 2128 3651 2156
rect 3635 2116 3651 2128
rect 3655 2116 3657 2156
rect 3669 2116 3671 2156
rect 3675 2116 3677 2156
rect 3733 2116 3735 2156
rect 3739 2136 3741 2156
rect 3753 2136 3755 2156
rect 3759 2136 3765 2156
rect 3769 2136 3773 2156
rect 3785 2136 3787 2156
rect 3791 2136 3797 2156
rect 3801 2136 3803 2156
rect 3815 2136 3819 2156
rect 3823 2136 3825 2156
rect 3863 2136 3865 2156
rect 3869 2136 3873 2156
rect 3877 2136 3879 2156
rect 3891 2136 3893 2156
rect 3897 2136 3903 2156
rect 3907 2136 3909 2156
rect 3921 2136 3925 2156
rect 3739 2116 3749 2136
rect 3912 2116 3925 2136
rect 3929 2116 3931 2156
rect 3969 2116 3971 2156
rect 3975 2136 3979 2156
rect 3991 2136 3993 2156
rect 3997 2136 4003 2156
rect 4007 2136 4009 2156
rect 4021 2136 4023 2156
rect 4027 2136 4031 2156
rect 4035 2136 4037 2156
rect 4075 2136 4077 2156
rect 4081 2136 4085 2156
rect 4097 2136 4099 2156
rect 4103 2136 4109 2156
rect 4113 2136 4115 2156
rect 4127 2136 4131 2156
rect 4135 2136 4141 2156
rect 4145 2136 4147 2156
rect 4159 2136 4161 2156
rect 3975 2116 3988 2136
rect 4151 2116 4161 2136
rect 4165 2116 4167 2156
rect 4244 2116 4246 2156
rect 4250 2116 4254 2156
rect 4258 2116 4260 2156
rect 4272 2116 4274 2156
rect 4278 2116 4282 2156
rect 4286 2116 4288 2156
rect 4329 2136 4331 2156
rect 4335 2136 4337 2156
rect 4403 2136 4405 2156
rect 4409 2136 4411 2156
rect 4423 2136 4425 2156
rect 4429 2136 4431 2156
rect 4483 2136 4485 2156
rect 4489 2136 4491 2156
rect 4503 2136 4505 2156
rect 4509 2136 4511 2156
rect 4549 2116 4551 2156
rect 4555 2136 4559 2156
rect 4571 2136 4573 2156
rect 4577 2136 4583 2156
rect 4587 2136 4589 2156
rect 4601 2136 4603 2156
rect 4607 2136 4611 2156
rect 4615 2136 4617 2156
rect 4655 2136 4657 2156
rect 4661 2136 4665 2156
rect 4677 2136 4679 2156
rect 4683 2136 4689 2156
rect 4693 2136 4695 2156
rect 4707 2136 4711 2156
rect 4715 2136 4721 2156
rect 4725 2136 4727 2156
rect 4739 2136 4741 2156
rect 4555 2116 4568 2136
rect 4731 2116 4741 2136
rect 4745 2116 4747 2156
rect 354 1762 368 1764
rect 64 1704 66 1744
rect 70 1704 74 1744
rect 78 1704 80 1744
rect 92 1704 94 1744
rect 98 1704 102 1744
rect 106 1704 108 1744
rect 149 1704 151 1744
rect 155 1732 171 1744
rect 155 1704 157 1732
rect 169 1704 171 1732
rect 175 1704 177 1744
rect 189 1704 191 1744
rect 195 1704 197 1744
rect 251 1704 253 1744
rect 257 1704 263 1744
rect 267 1704 269 1744
rect 366 1704 368 1762
rect 372 1704 376 1764
rect 380 1704 384 1764
rect 388 1704 390 1764
rect 432 1704 434 1744
rect 438 1704 442 1744
rect 446 1704 448 1744
rect 460 1704 462 1744
rect 466 1704 470 1744
rect 474 1704 476 1744
rect 549 1704 551 1744
rect 555 1704 561 1744
rect 565 1704 567 1744
rect 579 1704 581 1744
rect 585 1704 587 1744
rect 663 1704 665 1744
rect 669 1704 671 1744
rect 709 1704 711 1724
rect 715 1704 719 1724
rect 731 1704 733 1744
rect 737 1704 739 1744
rect 803 1704 805 1744
rect 809 1704 811 1744
rect 823 1704 825 1744
rect 829 1732 845 1744
rect 829 1704 831 1732
rect 843 1704 845 1732
rect 849 1704 851 1744
rect 889 1704 891 1744
rect 895 1732 911 1744
rect 895 1704 897 1732
rect 909 1704 911 1732
rect 915 1704 917 1744
rect 929 1704 931 1744
rect 935 1704 937 1744
rect 990 1704 992 1764
rect 996 1704 1000 1764
rect 1004 1704 1008 1764
rect 1012 1762 1026 1764
rect 1012 1704 1014 1762
rect 1089 1704 1091 1724
rect 1095 1704 1097 1724
rect 1150 1704 1152 1764
rect 1156 1704 1160 1764
rect 1164 1704 1168 1764
rect 1172 1762 1186 1764
rect 1172 1704 1174 1762
rect 1250 1704 1252 1764
rect 1256 1704 1260 1764
rect 1264 1704 1268 1764
rect 1272 1762 1286 1764
rect 1272 1704 1274 1762
rect 1363 1704 1365 1724
rect 1369 1704 1371 1724
rect 1444 1704 1446 1744
rect 1450 1704 1454 1744
rect 1458 1704 1460 1744
rect 1472 1704 1474 1744
rect 1478 1704 1482 1744
rect 1486 1704 1488 1744
rect 1530 1704 1532 1764
rect 1536 1704 1540 1764
rect 1544 1704 1548 1764
rect 1552 1762 1566 1764
rect 1552 1704 1554 1762
rect 1774 1762 1788 1764
rect 1629 1704 1631 1724
rect 1635 1704 1637 1724
rect 1703 1704 1705 1744
rect 1709 1704 1711 1744
rect 1786 1704 1788 1762
rect 1792 1704 1796 1764
rect 1800 1704 1804 1764
rect 1808 1704 1810 1764
rect 1849 1704 1851 1744
rect 1855 1704 1861 1744
rect 1865 1704 1867 1744
rect 1879 1704 1881 1744
rect 1885 1704 1887 1744
rect 1953 1704 1955 1744
rect 1959 1724 1969 1744
rect 2132 1724 2145 1744
rect 1959 1704 1961 1724
rect 1973 1704 1975 1724
rect 1979 1704 1985 1724
rect 1989 1704 1993 1724
rect 2005 1704 2007 1724
rect 2011 1704 2017 1724
rect 2021 1704 2023 1724
rect 2035 1704 2039 1724
rect 2043 1704 2045 1724
rect 2083 1704 2085 1724
rect 2089 1704 2093 1724
rect 2097 1704 2099 1724
rect 2111 1704 2113 1724
rect 2117 1704 2123 1724
rect 2127 1704 2129 1724
rect 2141 1704 2145 1724
rect 2149 1704 2151 1744
rect 2203 1704 2205 1724
rect 2209 1704 2211 1724
rect 2223 1704 2225 1724
rect 2229 1704 2231 1724
rect 2269 1704 2271 1724
rect 2275 1704 2277 1724
rect 2329 1704 2331 1744
rect 2335 1732 2351 1744
rect 2335 1704 2337 1732
rect 2349 1704 2351 1732
rect 2355 1704 2357 1744
rect 2369 1704 2371 1744
rect 2375 1704 2377 1744
rect 2429 1704 2431 1724
rect 2435 1704 2437 1724
rect 2449 1704 2451 1724
rect 2455 1704 2457 1724
rect 2509 1704 2511 1724
rect 2515 1704 2517 1724
rect 2529 1704 2531 1724
rect 2535 1704 2537 1724
rect 2589 1704 2591 1744
rect 2595 1732 2611 1744
rect 2595 1704 2597 1732
rect 2609 1704 2611 1732
rect 2615 1704 2617 1744
rect 2629 1704 2631 1744
rect 2635 1704 2637 1744
rect 2711 1704 2713 1744
rect 2717 1704 2723 1744
rect 2727 1704 2729 1744
rect 2783 1704 2785 1724
rect 2789 1704 2791 1724
rect 2803 1704 2805 1724
rect 2809 1704 2811 1724
rect 2849 1704 2851 1744
rect 2855 1732 2871 1744
rect 2855 1704 2857 1732
rect 2869 1704 2871 1732
rect 2875 1704 2877 1744
rect 2889 1704 2891 1744
rect 2895 1704 2897 1744
rect 2949 1704 2951 1724
rect 2955 1704 2957 1724
rect 3023 1704 3025 1724
rect 3029 1704 3031 1724
rect 3043 1704 3045 1724
rect 3049 1704 3051 1724
rect 3089 1704 3091 1744
rect 3095 1724 3108 1744
rect 3271 1724 3281 1744
rect 3095 1704 3099 1724
rect 3111 1704 3113 1724
rect 3117 1704 3123 1724
rect 3127 1704 3129 1724
rect 3141 1704 3143 1724
rect 3147 1704 3151 1724
rect 3155 1704 3157 1724
rect 3195 1704 3197 1724
rect 3201 1704 3205 1724
rect 3217 1704 3219 1724
rect 3223 1704 3229 1724
rect 3233 1704 3235 1724
rect 3247 1704 3251 1724
rect 3255 1704 3261 1724
rect 3265 1704 3267 1724
rect 3279 1704 3281 1724
rect 3285 1704 3287 1744
rect 3329 1704 3331 1744
rect 3335 1732 3351 1744
rect 3335 1704 3337 1732
rect 3349 1704 3351 1732
rect 3355 1704 3357 1744
rect 3369 1704 3371 1744
rect 3375 1704 3377 1744
rect 3431 1704 3433 1744
rect 3437 1704 3443 1744
rect 3447 1704 3449 1744
rect 3509 1704 3511 1744
rect 3515 1724 3528 1744
rect 3691 1724 3701 1744
rect 3515 1704 3519 1724
rect 3531 1704 3533 1724
rect 3537 1704 3543 1724
rect 3547 1704 3549 1724
rect 3561 1704 3563 1724
rect 3567 1704 3571 1724
rect 3575 1704 3577 1724
rect 3615 1704 3617 1724
rect 3621 1704 3625 1724
rect 3637 1704 3639 1724
rect 3643 1704 3649 1724
rect 3653 1704 3655 1724
rect 3667 1704 3671 1724
rect 3675 1704 3681 1724
rect 3685 1704 3687 1724
rect 3699 1704 3701 1724
rect 3705 1704 3707 1744
rect 3749 1704 3751 1724
rect 3755 1704 3759 1724
rect 3771 1704 3773 1744
rect 3777 1704 3779 1744
rect 3851 1704 3853 1744
rect 3857 1704 3863 1744
rect 3867 1704 3869 1744
rect 3923 1704 3925 1744
rect 3929 1704 3931 1744
rect 3943 1704 3945 1744
rect 3949 1732 3965 1744
rect 3949 1704 3951 1732
rect 3963 1704 3965 1732
rect 3969 1704 3971 1744
rect 4023 1704 4025 1744
rect 4029 1704 4031 1744
rect 4043 1704 4045 1744
rect 4049 1732 4065 1744
rect 4049 1704 4051 1732
rect 4063 1704 4065 1732
rect 4069 1704 4071 1744
rect 4139 1724 4151 1744
rect 4109 1704 4111 1724
rect 4115 1704 4117 1724
rect 4129 1704 4131 1724
rect 4135 1704 4137 1724
rect 4149 1704 4151 1724
rect 4155 1704 4157 1744
rect 4223 1704 4225 1724
rect 4229 1704 4231 1724
rect 4272 1704 4274 1744
rect 4278 1704 4282 1744
rect 4286 1704 4288 1744
rect 4300 1704 4304 1724
rect 4308 1704 4310 1724
rect 4383 1704 4385 1724
rect 4389 1704 4391 1724
rect 4403 1704 4405 1724
rect 4409 1704 4411 1724
rect 4449 1704 4451 1744
rect 4455 1724 4468 1744
rect 4631 1724 4641 1744
rect 4455 1704 4459 1724
rect 4471 1704 4473 1724
rect 4477 1704 4483 1724
rect 4487 1704 4489 1724
rect 4501 1704 4503 1724
rect 4507 1704 4511 1724
rect 4515 1704 4517 1724
rect 4555 1704 4557 1724
rect 4561 1704 4565 1724
rect 4577 1704 4579 1724
rect 4583 1704 4589 1724
rect 4593 1704 4595 1724
rect 4607 1704 4611 1724
rect 4615 1704 4621 1724
rect 4625 1704 4627 1724
rect 4639 1704 4641 1724
rect 4645 1704 4647 1744
rect 4711 1704 4713 1744
rect 4717 1704 4723 1744
rect 4727 1704 4729 1744
rect 43 1656 45 1676
rect 49 1656 51 1676
rect 110 1656 112 1676
rect 116 1656 120 1676
rect 132 1636 134 1676
rect 138 1636 142 1676
rect 146 1636 148 1676
rect 190 1616 192 1676
rect 196 1616 200 1676
rect 204 1616 208 1676
rect 212 1618 214 1676
rect 291 1636 293 1676
rect 297 1636 303 1676
rect 307 1636 309 1676
rect 383 1636 385 1676
rect 389 1636 391 1676
rect 403 1636 405 1676
rect 409 1648 411 1676
rect 423 1648 425 1676
rect 409 1636 425 1648
rect 429 1636 431 1676
rect 481 1636 483 1676
rect 487 1636 489 1676
rect 501 1656 505 1676
rect 509 1656 511 1676
rect 563 1656 565 1676
rect 569 1656 571 1676
rect 212 1616 226 1618
rect 610 1616 612 1676
rect 616 1616 620 1676
rect 624 1616 628 1676
rect 632 1618 634 1676
rect 712 1636 714 1676
rect 718 1636 722 1676
rect 726 1636 728 1676
rect 740 1656 744 1676
rect 748 1656 750 1676
rect 632 1616 646 1618
rect 810 1616 812 1676
rect 816 1616 820 1676
rect 824 1616 828 1676
rect 832 1618 834 1676
rect 912 1636 914 1676
rect 918 1636 922 1676
rect 926 1636 928 1676
rect 940 1656 944 1676
rect 948 1656 950 1676
rect 832 1616 846 1618
rect 1010 1616 1012 1676
rect 1016 1616 1020 1676
rect 1024 1616 1028 1676
rect 1032 1618 1034 1676
rect 1123 1636 1125 1676
rect 1129 1636 1131 1676
rect 1143 1636 1145 1676
rect 1149 1648 1151 1676
rect 1163 1648 1165 1676
rect 1149 1636 1165 1648
rect 1169 1636 1171 1676
rect 1032 1616 1046 1618
rect 1210 1616 1212 1676
rect 1216 1616 1220 1676
rect 1224 1616 1228 1676
rect 1232 1618 1234 1676
rect 1312 1636 1314 1676
rect 1318 1636 1322 1676
rect 1326 1636 1328 1676
rect 1340 1656 1344 1676
rect 1348 1656 1350 1676
rect 1423 1656 1425 1676
rect 1429 1656 1431 1676
rect 1232 1616 1246 1618
rect 1470 1616 1472 1676
rect 1476 1616 1480 1676
rect 1484 1616 1488 1676
rect 1492 1618 1494 1676
rect 1572 1636 1574 1676
rect 1578 1636 1582 1676
rect 1586 1636 1588 1676
rect 1600 1656 1604 1676
rect 1608 1656 1610 1676
rect 1492 1616 1506 1618
rect 1670 1616 1672 1676
rect 1676 1616 1680 1676
rect 1684 1616 1688 1676
rect 1692 1618 1694 1676
rect 1769 1636 1771 1676
rect 1775 1648 1777 1676
rect 1789 1648 1791 1676
rect 1775 1636 1791 1648
rect 1795 1636 1797 1676
rect 1809 1636 1811 1676
rect 1815 1636 1817 1676
rect 1890 1656 1892 1676
rect 1896 1656 1900 1676
rect 1692 1616 1706 1618
rect 1912 1636 1914 1676
rect 1918 1636 1922 1676
rect 1926 1636 1928 1676
rect 1969 1656 1971 1676
rect 1975 1656 1977 1676
rect 2030 1616 2032 1676
rect 2036 1616 2040 1676
rect 2044 1616 2048 1676
rect 2052 1618 2054 1676
rect 2143 1636 2145 1676
rect 2149 1636 2151 1676
rect 2163 1636 2165 1676
rect 2169 1648 2171 1676
rect 2183 1648 2185 1676
rect 2169 1636 2185 1648
rect 2189 1636 2191 1676
rect 2229 1656 2231 1676
rect 2235 1656 2237 1676
rect 2052 1616 2066 1618
rect 2289 1636 2291 1676
rect 2295 1656 2299 1676
rect 2311 1656 2313 1676
rect 2317 1656 2323 1676
rect 2327 1656 2329 1676
rect 2341 1656 2343 1676
rect 2347 1656 2351 1676
rect 2355 1656 2357 1676
rect 2395 1656 2397 1676
rect 2401 1656 2405 1676
rect 2417 1656 2419 1676
rect 2423 1656 2429 1676
rect 2433 1656 2435 1676
rect 2447 1656 2451 1676
rect 2455 1656 2461 1676
rect 2465 1656 2467 1676
rect 2479 1656 2481 1676
rect 2295 1636 2308 1656
rect 2471 1636 2481 1656
rect 2485 1636 2487 1676
rect 2543 1636 2545 1676
rect 2549 1636 2551 1676
rect 2563 1636 2565 1676
rect 2569 1648 2571 1676
rect 2583 1648 2585 1676
rect 2569 1636 2585 1648
rect 2589 1636 2591 1676
rect 2653 1636 2655 1676
rect 2659 1636 2661 1676
rect 2673 1636 2675 1676
rect 2679 1636 2685 1676
rect 2689 1636 2691 1676
rect 2729 1656 2731 1676
rect 2735 1656 2737 1676
rect 2749 1656 2751 1676
rect 2755 1656 2757 1676
rect 2812 1636 2814 1676
rect 2818 1636 2822 1676
rect 2826 1636 2828 1676
rect 2840 1656 2844 1676
rect 2848 1656 2850 1676
rect 2923 1656 2925 1676
rect 2929 1656 2931 1676
rect 2943 1656 2945 1676
rect 2949 1656 2951 1676
rect 3003 1656 3005 1676
rect 3009 1656 3011 1676
rect 3063 1656 3065 1676
rect 3069 1656 3071 1676
rect 3109 1636 3111 1676
rect 3115 1648 3117 1676
rect 3129 1648 3131 1676
rect 3115 1636 3131 1648
rect 3135 1636 3137 1676
rect 3149 1636 3151 1676
rect 3155 1636 3157 1676
rect 3211 1636 3213 1676
rect 3217 1636 3223 1676
rect 3227 1636 3229 1676
rect 3311 1636 3313 1676
rect 3317 1636 3323 1676
rect 3327 1636 3329 1676
rect 3383 1636 3385 1676
rect 3389 1636 3391 1676
rect 3403 1636 3405 1676
rect 3409 1648 3411 1676
rect 3423 1648 3425 1676
rect 3409 1636 3425 1648
rect 3429 1636 3431 1676
rect 3473 1636 3475 1676
rect 3479 1656 3481 1676
rect 3493 1656 3495 1676
rect 3499 1656 3505 1676
rect 3509 1656 3513 1676
rect 3525 1656 3527 1676
rect 3531 1656 3537 1676
rect 3541 1656 3543 1676
rect 3555 1656 3559 1676
rect 3563 1656 3565 1676
rect 3603 1656 3605 1676
rect 3609 1656 3613 1676
rect 3617 1656 3619 1676
rect 3631 1656 3633 1676
rect 3637 1656 3643 1676
rect 3647 1656 3649 1676
rect 3661 1656 3665 1676
rect 3479 1636 3489 1656
rect 3652 1636 3665 1656
rect 3669 1636 3671 1676
rect 3709 1656 3711 1676
rect 3715 1656 3717 1676
rect 3783 1656 3785 1676
rect 3789 1656 3791 1676
rect 3843 1636 3845 1676
rect 3849 1636 3851 1676
rect 3863 1636 3865 1676
rect 3869 1648 3871 1676
rect 3883 1648 3885 1676
rect 3869 1636 3885 1648
rect 3889 1636 3891 1676
rect 3929 1656 3931 1676
rect 3935 1656 3937 1676
rect 3949 1656 3951 1676
rect 3955 1656 3957 1676
rect 4009 1656 4011 1676
rect 4015 1656 4017 1676
rect 4029 1656 4031 1676
rect 4035 1656 4037 1676
rect 4089 1656 4091 1676
rect 4095 1656 4097 1676
rect 4152 1636 4154 1676
rect 4158 1636 4162 1676
rect 4166 1636 4168 1676
rect 4180 1656 4184 1676
rect 4188 1656 4190 1676
rect 4249 1656 4251 1676
rect 4255 1656 4257 1676
rect 4269 1656 4271 1676
rect 4275 1656 4277 1676
rect 4332 1636 4334 1676
rect 4338 1636 4342 1676
rect 4346 1636 4348 1676
rect 4360 1656 4364 1676
rect 4368 1656 4370 1676
rect 4429 1656 4431 1676
rect 4435 1656 4437 1676
rect 4489 1656 4491 1676
rect 4495 1656 4497 1676
rect 4563 1656 4565 1676
rect 4569 1656 4571 1676
rect 4609 1636 4611 1676
rect 4615 1648 4617 1676
rect 4629 1648 4631 1676
rect 4615 1636 4631 1648
rect 4635 1636 4637 1676
rect 4649 1636 4651 1676
rect 4655 1636 4657 1676
rect 4711 1636 4713 1676
rect 4717 1636 4723 1676
rect 4727 1636 4729 1676
rect 50 1224 52 1244
rect 56 1224 60 1244
rect 72 1224 74 1264
rect 78 1224 82 1264
rect 86 1224 88 1264
rect 130 1224 132 1284
rect 136 1224 140 1284
rect 144 1224 148 1284
rect 152 1282 166 1284
rect 152 1224 154 1282
rect 230 1224 232 1284
rect 236 1224 240 1284
rect 244 1224 248 1284
rect 252 1282 266 1284
rect 252 1224 254 1282
rect 351 1224 353 1264
rect 357 1224 363 1264
rect 367 1224 369 1264
rect 409 1224 411 1264
rect 415 1252 431 1264
rect 415 1224 417 1252
rect 429 1224 431 1252
rect 435 1224 437 1264
rect 449 1224 451 1264
rect 455 1224 457 1264
rect 512 1224 514 1264
rect 518 1224 522 1264
rect 526 1224 528 1264
rect 1094 1282 1108 1284
rect 540 1224 544 1244
rect 548 1224 550 1244
rect 609 1224 611 1264
rect 615 1252 631 1264
rect 615 1224 617 1252
rect 629 1224 631 1252
rect 635 1224 637 1264
rect 649 1224 651 1264
rect 655 1224 657 1264
rect 709 1224 711 1264
rect 715 1252 731 1264
rect 715 1224 717 1252
rect 729 1224 731 1252
rect 735 1224 737 1264
rect 749 1224 751 1264
rect 755 1224 757 1264
rect 809 1224 811 1264
rect 815 1224 821 1264
rect 825 1224 827 1264
rect 839 1224 841 1264
rect 845 1224 847 1264
rect 931 1224 933 1264
rect 937 1224 943 1264
rect 947 1224 949 1264
rect 991 1224 993 1264
rect 997 1224 1003 1264
rect 1007 1224 1009 1264
rect 1106 1224 1108 1282
rect 1112 1224 1116 1284
rect 1120 1224 1124 1284
rect 1128 1224 1130 1284
rect 1183 1224 1185 1244
rect 1189 1224 1191 1244
rect 1253 1224 1255 1264
rect 1259 1224 1261 1264
rect 1273 1224 1275 1264
rect 1279 1224 1285 1264
rect 1289 1224 1291 1264
rect 1329 1224 1331 1264
rect 1335 1252 1351 1264
rect 1335 1224 1337 1252
rect 1349 1224 1351 1252
rect 1355 1224 1357 1264
rect 1369 1224 1371 1264
rect 1375 1224 1377 1264
rect 1443 1224 1445 1264
rect 1449 1224 1451 1264
rect 1463 1224 1465 1264
rect 1469 1252 1485 1264
rect 1469 1224 1471 1252
rect 1483 1224 1485 1252
rect 1489 1224 1491 1264
rect 1531 1224 1533 1264
rect 1537 1224 1543 1264
rect 1547 1224 1549 1264
rect 1609 1224 1611 1264
rect 1615 1252 1631 1264
rect 1615 1224 1617 1252
rect 1629 1224 1631 1252
rect 1635 1224 1637 1264
rect 1649 1224 1651 1264
rect 1655 1224 1657 1264
rect 1711 1224 1713 1264
rect 1717 1224 1723 1264
rect 1727 1224 1729 1264
rect 1792 1224 1794 1264
rect 1798 1224 1802 1264
rect 1806 1224 1808 1264
rect 1820 1224 1824 1244
rect 1828 1224 1830 1244
rect 1890 1224 1892 1284
rect 1896 1224 1900 1284
rect 1904 1224 1908 1284
rect 1912 1282 1926 1284
rect 1912 1224 1914 1282
rect 1989 1224 1991 1264
rect 1995 1252 2011 1264
rect 1995 1224 1997 1252
rect 2009 1224 2011 1252
rect 2015 1224 2017 1264
rect 2029 1224 2031 1264
rect 2035 1224 2037 1264
rect 2089 1224 2091 1244
rect 2095 1224 2097 1244
rect 2150 1224 2152 1284
rect 2156 1224 2160 1284
rect 2164 1224 2168 1284
rect 2172 1282 2186 1284
rect 2172 1224 2174 1282
rect 2251 1224 2253 1264
rect 2257 1224 2263 1264
rect 2267 1224 2269 1264
rect 2359 1244 2371 1264
rect 2329 1224 2331 1244
rect 2335 1224 2337 1244
rect 2349 1224 2351 1244
rect 2355 1224 2357 1244
rect 2369 1224 2371 1244
rect 2375 1224 2377 1264
rect 2451 1224 2453 1264
rect 2457 1224 2463 1264
rect 2467 1224 2469 1264
rect 2509 1224 2511 1244
rect 2515 1224 2517 1244
rect 2581 1224 2583 1264
rect 2587 1224 2589 1264
rect 2601 1224 2605 1244
rect 2609 1224 2611 1244
rect 2649 1224 2651 1264
rect 2655 1252 2671 1264
rect 2655 1224 2657 1252
rect 2669 1224 2671 1252
rect 2675 1224 2677 1264
rect 2689 1224 2691 1264
rect 2695 1224 2697 1264
rect 2763 1224 2765 1264
rect 2769 1236 2771 1264
rect 2783 1236 2785 1264
rect 2769 1224 2785 1236
rect 2789 1224 2791 1264
rect 2803 1224 2805 1264
rect 2809 1254 2825 1264
rect 2809 1224 2811 1254
rect 2823 1224 2825 1254
rect 2829 1224 2831 1264
rect 2873 1224 2875 1264
rect 2879 1244 2889 1264
rect 3052 1244 3065 1264
rect 2879 1224 2881 1244
rect 2893 1224 2895 1244
rect 2899 1224 2905 1244
rect 2909 1224 2913 1244
rect 2925 1224 2927 1244
rect 2931 1224 2937 1244
rect 2941 1224 2943 1244
rect 2955 1224 2959 1244
rect 2963 1224 2965 1244
rect 3003 1224 3005 1244
rect 3009 1224 3013 1244
rect 3017 1224 3019 1244
rect 3031 1224 3033 1244
rect 3037 1224 3043 1244
rect 3047 1224 3049 1244
rect 3061 1224 3065 1244
rect 3069 1224 3071 1264
rect 3123 1224 3125 1244
rect 3129 1224 3131 1244
rect 3143 1224 3145 1244
rect 3149 1224 3151 1244
rect 3210 1224 3212 1244
rect 3216 1224 3220 1244
rect 3232 1224 3234 1264
rect 3238 1224 3242 1264
rect 3246 1224 3248 1264
rect 3293 1224 3295 1264
rect 3299 1244 3309 1264
rect 3472 1244 3485 1264
rect 3299 1224 3301 1244
rect 3313 1224 3315 1244
rect 3319 1224 3325 1244
rect 3329 1224 3333 1244
rect 3345 1224 3347 1244
rect 3351 1224 3357 1244
rect 3361 1224 3363 1244
rect 3375 1224 3379 1244
rect 3383 1224 3385 1244
rect 3423 1224 3425 1244
rect 3429 1224 3433 1244
rect 3437 1224 3439 1244
rect 3451 1224 3453 1244
rect 3457 1224 3463 1244
rect 3467 1224 3469 1244
rect 3481 1224 3485 1244
rect 3489 1224 3491 1264
rect 3543 1224 3545 1244
rect 3549 1224 3551 1244
rect 3603 1224 3605 1244
rect 3609 1224 3611 1244
rect 3623 1224 3625 1244
rect 3629 1224 3631 1244
rect 3683 1224 3685 1244
rect 3689 1224 3691 1244
rect 3703 1224 3705 1244
rect 3709 1224 3711 1244
rect 3749 1224 3751 1244
rect 3755 1224 3757 1244
rect 3809 1224 3811 1264
rect 3815 1244 3828 1264
rect 3991 1244 4001 1264
rect 3815 1224 3819 1244
rect 3831 1224 3833 1244
rect 3837 1224 3843 1244
rect 3847 1224 3849 1244
rect 3861 1224 3863 1244
rect 3867 1224 3871 1244
rect 3875 1224 3877 1244
rect 3915 1224 3917 1244
rect 3921 1224 3925 1244
rect 3937 1224 3939 1244
rect 3943 1224 3949 1244
rect 3953 1224 3955 1244
rect 3967 1224 3971 1244
rect 3975 1224 3981 1244
rect 3985 1224 3987 1244
rect 3999 1224 4001 1244
rect 4005 1224 4007 1264
rect 4049 1224 4051 1264
rect 4055 1252 4071 1264
rect 4055 1224 4057 1252
rect 4069 1224 4071 1252
rect 4075 1224 4077 1264
rect 4089 1224 4091 1264
rect 4095 1224 4097 1264
rect 4151 1224 4153 1264
rect 4157 1224 4163 1264
rect 4167 1224 4169 1264
rect 4241 1224 4243 1264
rect 4247 1224 4249 1264
rect 4261 1224 4265 1244
rect 4269 1224 4271 1244
rect 4331 1224 4333 1264
rect 4337 1224 4343 1264
rect 4347 1224 4349 1264
rect 4403 1224 4405 1264
rect 4409 1224 4411 1264
rect 4423 1224 4425 1264
rect 4429 1252 4445 1264
rect 4429 1224 4431 1252
rect 4443 1224 4445 1252
rect 4449 1224 4451 1264
rect 4503 1224 4505 1264
rect 4509 1224 4511 1264
rect 4523 1224 4525 1264
rect 4529 1252 4545 1264
rect 4529 1224 4531 1252
rect 4543 1224 4545 1252
rect 4549 1224 4551 1264
rect 4589 1224 4591 1244
rect 4595 1224 4597 1244
rect 4609 1224 4611 1244
rect 4615 1224 4617 1244
rect 4669 1224 4671 1244
rect 4675 1224 4677 1244
rect 4743 1224 4745 1244
rect 4749 1224 4751 1244
rect 43 1156 45 1196
rect 49 1156 51 1196
rect 63 1156 65 1196
rect 69 1168 71 1196
rect 83 1168 85 1196
rect 69 1156 85 1168
rect 89 1156 91 1196
rect 129 1156 131 1196
rect 135 1168 137 1196
rect 149 1168 151 1196
rect 135 1156 151 1168
rect 155 1156 157 1196
rect 169 1156 171 1196
rect 175 1156 177 1196
rect 230 1136 232 1196
rect 236 1136 240 1196
rect 244 1136 248 1196
rect 252 1138 254 1196
rect 332 1156 334 1196
rect 338 1156 342 1196
rect 346 1156 348 1196
rect 360 1176 364 1196
rect 368 1176 370 1196
rect 252 1136 266 1138
rect 430 1136 432 1196
rect 436 1136 440 1196
rect 444 1136 448 1196
rect 452 1138 454 1196
rect 532 1156 534 1196
rect 538 1156 542 1196
rect 546 1156 548 1196
rect 560 1176 564 1196
rect 568 1176 570 1196
rect 452 1136 466 1138
rect 651 1156 653 1196
rect 657 1156 663 1196
rect 667 1156 669 1196
rect 733 1156 735 1196
rect 739 1156 741 1196
rect 753 1156 755 1196
rect 759 1156 765 1196
rect 769 1156 771 1196
rect 846 1138 848 1196
rect 834 1136 848 1138
rect 852 1136 856 1196
rect 860 1136 864 1196
rect 868 1136 870 1196
rect 923 1156 925 1196
rect 929 1156 931 1196
rect 943 1156 945 1196
rect 949 1168 951 1196
rect 963 1168 965 1196
rect 949 1156 965 1168
rect 969 1156 971 1196
rect 1009 1156 1011 1196
rect 1015 1168 1017 1196
rect 1029 1168 1031 1196
rect 1015 1156 1031 1168
rect 1035 1156 1037 1196
rect 1049 1156 1051 1196
rect 1055 1156 1057 1196
rect 1123 1156 1125 1196
rect 1129 1156 1131 1196
rect 1143 1156 1145 1196
rect 1149 1168 1151 1196
rect 1163 1168 1165 1196
rect 1149 1156 1165 1168
rect 1169 1156 1171 1196
rect 1231 1156 1233 1196
rect 1237 1156 1243 1196
rect 1247 1156 1249 1196
rect 1313 1156 1315 1196
rect 1319 1156 1321 1196
rect 1333 1156 1335 1196
rect 1339 1156 1345 1196
rect 1349 1156 1351 1196
rect 1391 1156 1393 1196
rect 1397 1156 1403 1196
rect 1407 1156 1409 1196
rect 1483 1156 1485 1196
rect 1489 1156 1491 1196
rect 1551 1156 1553 1196
rect 1557 1156 1563 1196
rect 1567 1156 1569 1196
rect 1631 1156 1633 1196
rect 1637 1156 1643 1196
rect 1647 1156 1649 1196
rect 1690 1136 1692 1196
rect 1696 1136 1700 1196
rect 1704 1136 1708 1196
rect 1712 1138 1714 1196
rect 1811 1156 1813 1196
rect 1817 1156 1823 1196
rect 1827 1156 1829 1196
rect 1712 1136 1726 1138
rect 1870 1136 1872 1196
rect 1876 1136 1880 1196
rect 1884 1136 1888 1196
rect 1892 1138 1894 1196
rect 1971 1156 1973 1196
rect 1977 1156 1983 1196
rect 1987 1156 1989 1196
rect 2084 1156 2086 1196
rect 2090 1156 2094 1196
rect 2098 1156 2100 1196
rect 2112 1156 2114 1196
rect 2118 1156 2122 1196
rect 2126 1156 2128 1196
rect 1892 1136 1906 1138
rect 2206 1138 2208 1196
rect 2194 1136 2208 1138
rect 2212 1136 2216 1196
rect 2220 1136 2224 1196
rect 2228 1136 2230 1196
rect 2291 1156 2293 1196
rect 2297 1156 2303 1196
rect 2307 1156 2309 1196
rect 2352 1156 2354 1196
rect 2358 1156 2362 1196
rect 2366 1156 2368 1196
rect 2380 1176 2384 1196
rect 2388 1176 2390 1196
rect 2463 1176 2465 1196
rect 2469 1176 2471 1196
rect 2531 1156 2533 1196
rect 2537 1156 2543 1196
rect 2547 1156 2549 1196
rect 2603 1156 2605 1196
rect 2609 1184 2625 1196
rect 2609 1156 2611 1184
rect 2623 1156 2625 1184
rect 2629 1156 2631 1196
rect 2643 1156 2645 1196
rect 2649 1166 2651 1196
rect 2663 1166 2665 1196
rect 2649 1156 2665 1166
rect 2669 1156 2671 1196
rect 2709 1176 2711 1196
rect 2715 1176 2719 1196
rect 2731 1156 2733 1196
rect 2737 1156 2739 1196
rect 2793 1156 2795 1196
rect 2799 1176 2801 1196
rect 2813 1176 2815 1196
rect 2819 1176 2825 1196
rect 2829 1176 2833 1196
rect 2845 1176 2847 1196
rect 2851 1176 2857 1196
rect 2861 1176 2863 1196
rect 2875 1176 2879 1196
rect 2883 1176 2885 1196
rect 2923 1176 2925 1196
rect 2929 1176 2933 1196
rect 2937 1176 2939 1196
rect 2951 1176 2953 1196
rect 2957 1176 2963 1196
rect 2967 1176 2969 1196
rect 2981 1176 2985 1196
rect 2799 1156 2809 1176
rect 2972 1156 2985 1176
rect 2989 1156 2991 1196
rect 3031 1156 3033 1196
rect 3037 1156 3043 1196
rect 3047 1156 3049 1196
rect 3123 1156 3125 1196
rect 3129 1156 3131 1196
rect 3143 1156 3145 1196
rect 3149 1168 3151 1196
rect 3163 1168 3165 1196
rect 3149 1156 3165 1168
rect 3169 1156 3171 1196
rect 3209 1156 3211 1196
rect 3215 1156 3217 1196
rect 3229 1156 3231 1196
rect 3235 1156 3237 1196
rect 3249 1156 3251 1196
rect 3255 1156 3257 1196
rect 3269 1156 3271 1196
rect 3275 1156 3277 1196
rect 3341 1156 3343 1196
rect 3347 1156 3349 1196
rect 3361 1176 3365 1196
rect 3369 1176 3371 1196
rect 3409 1176 3411 1196
rect 3415 1176 3419 1196
rect 3431 1156 3433 1196
rect 3437 1156 3439 1196
rect 3489 1156 3491 1196
rect 3495 1156 3497 1196
rect 3509 1156 3511 1196
rect 3515 1156 3517 1196
rect 3529 1156 3531 1196
rect 3535 1156 3537 1196
rect 3549 1156 3551 1196
rect 3555 1156 3557 1196
rect 3569 1156 3571 1196
rect 3575 1156 3577 1196
rect 3589 1156 3591 1196
rect 3595 1156 3597 1196
rect 3609 1156 3611 1196
rect 3615 1156 3617 1196
rect 3629 1156 3631 1196
rect 3635 1156 3637 1196
rect 3689 1156 3691 1196
rect 3695 1156 3697 1196
rect 3709 1156 3711 1196
rect 3715 1156 3717 1196
rect 3729 1156 3731 1196
rect 3735 1156 3737 1196
rect 3749 1156 3751 1196
rect 3755 1156 3757 1196
rect 3769 1156 3771 1196
rect 3775 1156 3777 1196
rect 3789 1156 3791 1196
rect 3795 1156 3797 1196
rect 3809 1156 3811 1196
rect 3815 1156 3817 1196
rect 3829 1156 3831 1196
rect 3835 1156 3837 1196
rect 3889 1176 3891 1196
rect 3895 1176 3899 1196
rect 3911 1156 3913 1196
rect 3917 1156 3919 1196
rect 3971 1156 3973 1196
rect 3977 1156 3983 1196
rect 3987 1156 3989 1196
rect 4049 1156 4051 1196
rect 4055 1176 4059 1196
rect 4071 1176 4073 1196
rect 4077 1176 4083 1196
rect 4087 1176 4089 1196
rect 4101 1176 4103 1196
rect 4107 1176 4111 1196
rect 4115 1176 4117 1196
rect 4155 1176 4157 1196
rect 4161 1176 4165 1196
rect 4177 1176 4179 1196
rect 4183 1176 4189 1196
rect 4193 1176 4195 1196
rect 4207 1176 4211 1196
rect 4215 1176 4221 1196
rect 4225 1176 4227 1196
rect 4239 1176 4241 1196
rect 4055 1156 4068 1176
rect 4231 1156 4241 1176
rect 4245 1156 4247 1196
rect 4291 1156 4293 1196
rect 4297 1156 4303 1196
rect 4307 1156 4309 1196
rect 4369 1156 4371 1196
rect 4375 1168 4377 1196
rect 4389 1168 4391 1196
rect 4375 1156 4391 1168
rect 4395 1156 4397 1196
rect 4409 1156 4411 1196
rect 4415 1156 4417 1196
rect 4491 1156 4493 1196
rect 4497 1156 4503 1196
rect 4507 1156 4509 1196
rect 4549 1156 4551 1196
rect 4555 1168 4557 1196
rect 4569 1168 4571 1196
rect 4555 1156 4571 1168
rect 4575 1156 4577 1196
rect 4589 1156 4591 1196
rect 4595 1156 4597 1196
rect 4650 1136 4652 1196
rect 4656 1136 4660 1196
rect 4664 1136 4668 1196
rect 4672 1138 4674 1196
rect 4672 1136 4686 1138
rect 51 744 53 784
rect 57 744 63 784
rect 67 744 69 784
rect 133 744 135 784
rect 139 744 141 784
rect 153 744 155 784
rect 159 744 165 784
rect 169 744 171 784
rect 223 744 225 784
rect 229 744 231 784
rect 243 744 245 784
rect 249 772 265 784
rect 249 744 251 772
rect 263 744 265 772
rect 269 744 271 784
rect 344 744 346 784
rect 350 744 354 784
rect 358 744 360 784
rect 372 744 374 784
rect 378 744 382 784
rect 386 744 388 784
rect 441 744 443 784
rect 447 744 449 784
rect 461 744 465 764
rect 469 744 471 764
rect 509 744 511 764
rect 515 744 517 764
rect 583 744 585 764
rect 589 744 591 764
rect 650 744 652 764
rect 656 744 660 764
rect 672 744 674 784
rect 678 744 682 784
rect 686 744 688 784
rect 730 744 732 804
rect 736 744 740 804
rect 744 744 748 804
rect 752 802 766 804
rect 752 744 754 802
rect 1034 802 1048 804
rect 853 744 855 784
rect 859 744 861 784
rect 873 744 875 784
rect 879 744 885 784
rect 889 744 891 784
rect 931 744 933 784
rect 937 744 943 784
rect 947 744 949 784
rect 1046 744 1048 802
rect 1052 744 1056 804
rect 1060 744 1064 804
rect 1068 744 1070 804
rect 1234 802 1248 804
rect 1109 744 1111 784
rect 1115 772 1131 784
rect 1115 744 1117 772
rect 1129 744 1131 772
rect 1135 744 1137 784
rect 1149 744 1151 784
rect 1155 744 1157 784
rect 1246 744 1248 802
rect 1252 744 1256 804
rect 1260 744 1264 804
rect 1268 744 1270 804
rect 1309 744 1311 764
rect 1315 744 1317 764
rect 1369 744 1371 784
rect 1375 772 1391 784
rect 1375 744 1377 772
rect 1389 744 1391 772
rect 1395 744 1397 784
rect 1409 744 1411 784
rect 1415 744 1417 784
rect 1491 744 1493 784
rect 1497 744 1503 784
rect 1507 744 1509 784
rect 1551 744 1553 784
rect 1557 744 1563 784
rect 1567 744 1569 784
rect 1643 744 1645 784
rect 1649 744 1651 784
rect 1663 744 1665 784
rect 1669 772 1685 784
rect 1669 744 1671 772
rect 1683 744 1685 772
rect 1689 744 1691 784
rect 1729 744 1731 784
rect 1735 744 1741 784
rect 1745 744 1747 784
rect 1759 744 1761 784
rect 1765 744 1767 784
rect 1843 744 1845 764
rect 1849 744 1851 764
rect 1911 744 1913 784
rect 1917 744 1923 784
rect 1927 744 1929 784
rect 2054 802 2068 804
rect 1969 744 1971 764
rect 1975 744 1977 764
rect 2066 744 2068 802
rect 2072 744 2076 804
rect 2080 744 2084 804
rect 2088 744 2090 804
rect 2129 744 2131 764
rect 2135 744 2137 764
rect 2189 744 2191 784
rect 2195 772 2211 784
rect 2195 744 2197 772
rect 2209 744 2211 772
rect 2215 744 2217 784
rect 2229 744 2231 784
rect 2235 744 2237 784
rect 2310 744 2312 764
rect 2316 744 2320 764
rect 2332 744 2334 784
rect 2338 744 2342 784
rect 2346 744 2348 784
rect 2389 744 2391 764
rect 2395 744 2397 764
rect 2450 744 2452 804
rect 2456 744 2460 804
rect 2464 744 2468 804
rect 2472 802 2486 804
rect 2472 744 2474 802
rect 2574 802 2588 804
rect 2586 744 2588 802
rect 2592 744 2596 804
rect 2600 744 2604 804
rect 2608 744 2610 804
rect 2652 744 2654 784
rect 2658 744 2662 784
rect 2666 744 2668 784
rect 2680 744 2684 764
rect 2688 744 2690 764
rect 2771 744 2773 784
rect 2777 744 2783 784
rect 2787 744 2789 784
rect 2843 744 2845 784
rect 2849 756 2851 784
rect 2863 756 2865 784
rect 2849 744 2865 756
rect 2869 744 2871 784
rect 2883 744 2885 784
rect 2889 774 2905 784
rect 2889 744 2891 774
rect 2903 744 2905 774
rect 2909 744 2911 784
rect 2963 744 2965 764
rect 2969 744 2971 764
rect 3023 744 3025 764
rect 3029 744 3031 764
rect 3043 744 3045 764
rect 3049 744 3051 764
rect 3103 744 3105 764
rect 3109 744 3111 764
rect 3123 744 3125 764
rect 3129 744 3131 764
rect 3169 744 3171 764
rect 3175 744 3177 764
rect 3229 744 3231 784
rect 3235 772 3251 784
rect 3235 744 3237 772
rect 3249 744 3251 772
rect 3255 744 3257 784
rect 3269 744 3271 784
rect 3275 744 3277 784
rect 3331 744 3333 784
rect 3337 744 3343 784
rect 3347 744 3349 784
rect 3409 744 3411 784
rect 3415 764 3428 784
rect 3591 764 3601 784
rect 3415 744 3419 764
rect 3431 744 3433 764
rect 3437 744 3443 764
rect 3447 744 3449 764
rect 3461 744 3463 764
rect 3467 744 3471 764
rect 3475 744 3477 764
rect 3515 744 3517 764
rect 3521 744 3525 764
rect 3537 744 3539 764
rect 3543 744 3549 764
rect 3553 744 3555 764
rect 3567 744 3571 764
rect 3575 744 3581 764
rect 3585 744 3587 764
rect 3599 744 3601 764
rect 3605 744 3607 784
rect 3649 744 3651 764
rect 3655 744 3659 764
rect 3671 744 3673 784
rect 3677 744 3679 784
rect 3733 744 3735 784
rect 3739 764 3749 784
rect 3912 764 3925 784
rect 3739 744 3741 764
rect 3753 744 3755 764
rect 3759 744 3765 764
rect 3769 744 3773 764
rect 3785 744 3787 764
rect 3791 744 3797 764
rect 3801 744 3803 764
rect 3815 744 3819 764
rect 3823 744 3825 764
rect 3863 744 3865 764
rect 3869 744 3873 764
rect 3877 744 3879 764
rect 3891 744 3893 764
rect 3897 744 3903 764
rect 3907 744 3909 764
rect 3921 744 3925 764
rect 3929 744 3931 784
rect 3983 744 3985 784
rect 3989 744 3991 784
rect 4003 744 4005 784
rect 4009 772 4025 784
rect 4009 744 4011 772
rect 4023 744 4025 772
rect 4029 744 4031 784
rect 4069 744 4071 784
rect 4075 764 4088 784
rect 4251 764 4261 784
rect 4075 744 4079 764
rect 4091 744 4093 764
rect 4097 744 4103 764
rect 4107 744 4109 764
rect 4121 744 4123 764
rect 4127 744 4131 764
rect 4135 744 4137 764
rect 4175 744 4177 764
rect 4181 744 4185 764
rect 4197 744 4199 764
rect 4203 744 4209 764
rect 4213 744 4215 764
rect 4227 744 4231 764
rect 4235 744 4241 764
rect 4245 744 4247 764
rect 4259 744 4261 764
rect 4265 744 4267 784
rect 4313 744 4315 784
rect 4319 764 4329 784
rect 4492 764 4505 784
rect 4319 744 4321 764
rect 4333 744 4335 764
rect 4339 744 4345 764
rect 4349 744 4353 764
rect 4365 744 4367 764
rect 4371 744 4377 764
rect 4381 744 4383 764
rect 4395 744 4399 764
rect 4403 744 4405 764
rect 4443 744 4445 764
rect 4449 744 4453 764
rect 4457 744 4459 764
rect 4471 744 4473 764
rect 4477 744 4483 764
rect 4487 744 4489 764
rect 4501 744 4505 764
rect 4509 744 4511 784
rect 4549 744 4551 784
rect 4555 772 4571 784
rect 4555 744 4557 772
rect 4569 744 4571 772
rect 4575 744 4577 784
rect 4589 744 4591 784
rect 4595 744 4597 784
rect 4649 744 4651 784
rect 4655 772 4671 784
rect 4655 744 4657 772
rect 4669 744 4671 772
rect 4675 744 4677 784
rect 4689 744 4691 784
rect 4695 744 4697 784
rect 43 696 45 716
rect 49 696 51 716
rect 63 696 65 716
rect 69 696 71 716
rect 130 696 132 716
rect 136 696 140 716
rect 152 676 154 716
rect 158 676 162 716
rect 166 676 168 716
rect 209 696 211 716
rect 215 696 217 716
rect 290 696 292 716
rect 296 696 300 716
rect 312 676 314 716
rect 318 676 322 716
rect 326 676 328 716
rect 370 656 372 716
rect 376 656 380 716
rect 384 656 388 716
rect 392 658 394 716
rect 483 676 485 716
rect 489 676 491 716
rect 503 676 505 716
rect 509 688 511 716
rect 523 688 525 716
rect 509 676 525 688
rect 529 676 531 716
rect 581 676 583 716
rect 587 676 589 716
rect 601 696 605 716
rect 609 696 611 716
rect 392 656 406 658
rect 663 676 665 716
rect 669 676 671 716
rect 683 676 685 716
rect 689 688 691 716
rect 703 688 705 716
rect 689 676 705 688
rect 709 676 711 716
rect 761 676 763 716
rect 767 676 769 716
rect 781 696 785 716
rect 789 696 791 716
rect 829 676 831 716
rect 835 676 841 716
rect 845 676 847 716
rect 859 676 861 716
rect 865 676 867 716
rect 929 676 931 716
rect 935 688 937 716
rect 949 688 951 716
rect 935 676 951 688
rect 955 676 957 716
rect 969 676 971 716
rect 975 676 977 716
rect 1043 676 1045 716
rect 1049 676 1051 716
rect 1063 676 1065 716
rect 1069 688 1071 716
rect 1083 688 1085 716
rect 1069 676 1085 688
rect 1089 676 1091 716
rect 1143 676 1145 716
rect 1149 676 1151 716
rect 1192 676 1194 716
rect 1198 676 1202 716
rect 1206 676 1208 716
rect 1220 696 1224 716
rect 1228 696 1230 716
rect 1303 696 1305 716
rect 1309 696 1311 716
rect 1349 676 1351 716
rect 1355 688 1357 716
rect 1369 688 1371 716
rect 1355 676 1371 688
rect 1375 676 1377 716
rect 1389 676 1391 716
rect 1395 676 1397 716
rect 1449 676 1451 716
rect 1455 688 1457 716
rect 1469 688 1471 716
rect 1455 676 1471 688
rect 1475 676 1477 716
rect 1489 676 1491 716
rect 1495 676 1497 716
rect 1570 696 1572 716
rect 1576 696 1580 716
rect 1592 676 1594 716
rect 1598 676 1602 716
rect 1606 676 1608 716
rect 1652 676 1654 716
rect 1658 676 1662 716
rect 1666 676 1668 716
rect 1680 696 1684 716
rect 1688 696 1690 716
rect 1750 656 1752 716
rect 1756 656 1760 716
rect 1764 656 1768 716
rect 1772 658 1774 716
rect 1849 676 1851 716
rect 1855 688 1857 716
rect 1869 688 1871 716
rect 1855 676 1871 688
rect 1875 676 1877 716
rect 1889 676 1891 716
rect 1895 676 1897 716
rect 1970 696 1972 716
rect 1976 696 1980 716
rect 1772 656 1786 658
rect 1992 676 1994 716
rect 1998 676 2002 716
rect 2006 676 2008 716
rect 2049 676 2051 716
rect 2055 688 2057 716
rect 2069 688 2071 716
rect 2055 676 2071 688
rect 2075 676 2077 716
rect 2089 676 2091 716
rect 2095 676 2097 716
rect 2186 658 2188 716
rect 2174 656 2188 658
rect 2192 656 2196 716
rect 2200 656 2204 716
rect 2208 656 2210 716
rect 2263 676 2265 716
rect 2269 676 2271 716
rect 2283 676 2285 716
rect 2289 688 2291 716
rect 2303 688 2305 716
rect 2289 676 2305 688
rect 2309 676 2311 716
rect 2349 676 2351 716
rect 2355 688 2357 716
rect 2369 688 2371 716
rect 2355 676 2371 688
rect 2375 676 2377 716
rect 2389 676 2391 716
rect 2395 676 2397 716
rect 2450 656 2452 716
rect 2456 656 2460 716
rect 2464 656 2468 716
rect 2472 658 2474 716
rect 2472 656 2486 658
rect 2550 656 2552 716
rect 2556 656 2560 716
rect 2564 656 2568 716
rect 2572 658 2574 716
rect 2663 696 2665 716
rect 2669 696 2671 716
rect 2572 656 2586 658
rect 2710 656 2712 716
rect 2716 656 2720 716
rect 2724 656 2728 716
rect 2732 658 2734 716
rect 2813 676 2815 716
rect 2819 696 2821 716
rect 2833 696 2835 716
rect 2839 696 2845 716
rect 2849 696 2853 716
rect 2865 696 2867 716
rect 2871 696 2877 716
rect 2881 696 2883 716
rect 2895 696 2899 716
rect 2903 696 2905 716
rect 2943 696 2945 716
rect 2949 696 2953 716
rect 2957 696 2959 716
rect 2971 696 2973 716
rect 2977 696 2983 716
rect 2987 696 2989 716
rect 3001 696 3005 716
rect 2819 676 2829 696
rect 2732 656 2746 658
rect 2992 676 3005 696
rect 3009 676 3011 716
rect 3049 676 3051 716
rect 3055 688 3057 716
rect 3069 688 3071 716
rect 3055 676 3071 688
rect 3075 676 3077 716
rect 3089 676 3091 716
rect 3095 676 3097 716
rect 3149 696 3151 716
rect 3155 696 3157 716
rect 3209 696 3211 716
rect 3215 696 3217 716
rect 3270 656 3272 716
rect 3276 656 3280 716
rect 3284 656 3288 716
rect 3292 658 3294 716
rect 3383 696 3385 716
rect 3389 696 3391 716
rect 3292 656 3306 658
rect 3451 676 3453 716
rect 3457 676 3463 716
rect 3467 676 3469 716
rect 3523 676 3525 716
rect 3529 676 3531 716
rect 3543 676 3545 716
rect 3549 688 3551 716
rect 3563 688 3565 716
rect 3549 676 3565 688
rect 3569 676 3571 716
rect 3613 676 3615 716
rect 3619 696 3621 716
rect 3633 696 3635 716
rect 3639 696 3645 716
rect 3649 696 3653 716
rect 3665 696 3667 716
rect 3671 696 3677 716
rect 3681 696 3683 716
rect 3695 696 3699 716
rect 3703 696 3705 716
rect 3743 696 3745 716
rect 3749 696 3753 716
rect 3757 696 3759 716
rect 3771 696 3773 716
rect 3777 696 3783 716
rect 3787 696 3789 716
rect 3801 696 3805 716
rect 3619 676 3629 696
rect 3792 676 3805 696
rect 3809 676 3811 716
rect 3849 676 3851 716
rect 3855 688 3857 716
rect 3869 688 3871 716
rect 3855 676 3871 688
rect 3875 676 3877 716
rect 3889 676 3891 716
rect 3895 676 3897 716
rect 3971 676 3973 716
rect 3977 676 3983 716
rect 3987 676 3989 716
rect 4029 676 4031 716
rect 4035 696 4039 716
rect 4051 696 4053 716
rect 4057 696 4063 716
rect 4067 696 4069 716
rect 4081 696 4083 716
rect 4087 696 4091 716
rect 4095 696 4097 716
rect 4135 696 4137 716
rect 4141 696 4145 716
rect 4157 696 4159 716
rect 4163 696 4169 716
rect 4173 696 4175 716
rect 4187 696 4191 716
rect 4195 696 4201 716
rect 4205 696 4207 716
rect 4219 696 4221 716
rect 4035 676 4048 696
rect 4211 676 4221 696
rect 4225 676 4227 716
rect 4271 676 4273 716
rect 4277 676 4283 716
rect 4287 676 4289 716
rect 4351 676 4353 716
rect 4357 676 4363 716
rect 4367 676 4369 716
rect 4443 676 4445 716
rect 4449 676 4451 716
rect 4463 676 4465 716
rect 4469 688 4471 716
rect 4483 688 4485 716
rect 4469 676 4485 688
rect 4489 676 4491 716
rect 4533 676 4535 716
rect 4539 696 4541 716
rect 4553 696 4555 716
rect 4559 696 4565 716
rect 4569 696 4573 716
rect 4585 696 4587 716
rect 4591 696 4597 716
rect 4601 696 4603 716
rect 4615 696 4619 716
rect 4623 696 4625 716
rect 4663 696 4665 716
rect 4669 696 4673 716
rect 4677 696 4679 716
rect 4691 696 4693 716
rect 4697 696 4703 716
rect 4707 696 4709 716
rect 4721 696 4725 716
rect 4539 676 4549 696
rect 4712 676 4725 696
rect 4729 676 4731 716
rect 554 322 568 324
rect 31 264 33 304
rect 37 264 43 304
rect 47 264 49 304
rect 111 264 113 304
rect 117 264 123 304
rect 127 264 129 304
rect 211 264 213 304
rect 217 264 223 304
rect 227 264 229 304
rect 291 264 293 304
rect 297 264 303 304
rect 307 264 309 304
rect 373 264 375 304
rect 379 264 381 304
rect 393 264 395 304
rect 399 264 405 304
rect 409 264 411 304
rect 471 264 473 304
rect 477 264 483 304
rect 487 264 489 304
rect 566 264 568 322
rect 572 264 576 324
rect 580 264 584 324
rect 588 264 590 324
rect 664 264 666 304
rect 670 264 674 304
rect 678 264 680 304
rect 692 264 694 304
rect 698 264 702 304
rect 706 264 708 304
rect 763 264 765 284
rect 769 264 771 284
rect 783 264 785 284
rect 789 264 791 284
rect 851 264 853 304
rect 857 264 863 304
rect 867 264 869 304
rect 911 264 913 304
rect 917 264 923 304
rect 927 264 929 304
rect 1011 264 1013 304
rect 1017 264 1023 304
rect 1027 264 1029 304
rect 1091 264 1093 304
rect 1097 264 1103 304
rect 1107 264 1109 304
rect 1184 264 1186 304
rect 1190 264 1194 304
rect 1198 264 1200 304
rect 1212 264 1214 304
rect 1218 264 1222 304
rect 1226 264 1228 304
rect 1269 264 1271 304
rect 1275 292 1291 304
rect 1275 264 1277 292
rect 1289 264 1291 292
rect 1295 264 1297 304
rect 1309 264 1311 304
rect 1315 264 1317 304
rect 1383 264 1385 284
rect 1389 264 1391 284
rect 1403 264 1405 284
rect 1409 264 1411 284
rect 1449 264 1451 304
rect 1455 292 1471 304
rect 1455 264 1457 292
rect 1469 264 1471 292
rect 1475 264 1477 304
rect 1489 264 1491 304
rect 1495 264 1497 304
rect 1549 264 1551 284
rect 1555 264 1557 284
rect 1630 264 1632 284
rect 1636 264 1640 284
rect 1652 264 1654 304
rect 1658 264 1662 304
rect 1666 264 1668 304
rect 1709 264 1711 284
rect 1715 264 1717 284
rect 1770 264 1772 324
rect 1776 264 1780 324
rect 1784 264 1788 324
rect 1792 322 1806 324
rect 1792 264 1794 322
rect 1872 264 1874 304
rect 1878 264 1882 304
rect 1886 264 1888 304
rect 1900 264 1904 284
rect 1908 264 1910 284
rect 1971 264 1973 304
rect 1977 264 1983 304
rect 1987 264 1989 304
rect 2051 264 2053 304
rect 2057 264 2063 304
rect 2067 264 2069 304
rect 2131 264 2133 304
rect 2137 264 2143 304
rect 2147 264 2149 304
rect 2223 264 2225 284
rect 2229 264 2231 284
rect 2243 264 2245 284
rect 2249 264 2251 284
rect 2311 264 2313 304
rect 2317 264 2323 304
rect 2327 264 2329 304
rect 2369 264 2371 284
rect 2375 264 2377 284
rect 2389 264 2391 284
rect 2395 264 2397 284
rect 2450 264 2452 324
rect 2456 264 2460 324
rect 2464 264 2468 324
rect 2472 322 2486 324
rect 2472 264 2474 322
rect 2634 322 2648 324
rect 2563 264 2565 284
rect 2569 264 2571 284
rect 2646 264 2648 322
rect 2652 264 2656 324
rect 2660 264 2664 324
rect 2668 264 2670 324
rect 2712 264 2714 304
rect 2718 264 2722 304
rect 2726 264 2728 304
rect 2740 264 2744 284
rect 2748 264 2750 284
rect 2809 264 2811 284
rect 2815 264 2817 284
rect 2829 264 2831 284
rect 2835 264 2837 284
rect 2911 264 2913 304
rect 2917 264 2923 304
rect 2927 264 2929 304
rect 2983 264 2985 304
rect 2989 264 2991 304
rect 3003 264 3005 304
rect 3009 292 3025 304
rect 3009 264 3011 292
rect 3023 264 3025 292
rect 3029 264 3031 304
rect 3083 264 3085 304
rect 3089 264 3091 304
rect 3103 264 3105 304
rect 3109 292 3125 304
rect 3109 264 3111 292
rect 3123 264 3125 292
rect 3129 264 3131 304
rect 3183 264 3185 284
rect 3189 264 3191 284
rect 3203 264 3205 284
rect 3209 264 3211 284
rect 3263 264 3265 284
rect 3269 264 3271 284
rect 3323 264 3325 304
rect 3329 264 3331 304
rect 3343 264 3345 304
rect 3349 292 3365 304
rect 3349 264 3351 292
rect 3363 264 3365 292
rect 3369 264 3371 304
rect 3430 264 3432 284
rect 3436 264 3440 284
rect 3452 264 3454 304
rect 3458 264 3462 304
rect 3466 264 3468 304
rect 3619 284 3631 304
rect 3523 264 3525 284
rect 3529 264 3531 284
rect 3543 264 3545 284
rect 3549 264 3551 284
rect 3589 264 3591 284
rect 3595 264 3597 284
rect 3609 264 3611 284
rect 3615 264 3617 284
rect 3629 264 3631 284
rect 3635 264 3637 304
rect 3691 264 3693 304
rect 3697 264 3703 304
rect 3707 264 3709 304
rect 3771 264 3773 304
rect 3777 264 3783 304
rect 3787 264 3789 304
rect 3863 264 3865 304
rect 3869 264 3871 304
rect 3883 264 3885 304
rect 3889 292 3905 304
rect 3889 264 3891 292
rect 3903 264 3905 292
rect 3909 264 3911 304
rect 3963 264 3965 284
rect 3969 264 3971 284
rect 4023 264 4025 284
rect 4029 264 4031 284
rect 4069 264 4071 304
rect 4075 284 4088 304
rect 4251 284 4261 304
rect 4075 264 4079 284
rect 4091 264 4093 284
rect 4097 264 4103 284
rect 4107 264 4109 284
rect 4121 264 4123 284
rect 4127 264 4131 284
rect 4135 264 4137 284
rect 4175 264 4177 284
rect 4181 264 4185 284
rect 4197 264 4199 284
rect 4203 264 4209 284
rect 4213 264 4215 284
rect 4227 264 4231 284
rect 4235 264 4241 284
rect 4245 264 4247 284
rect 4259 264 4261 284
rect 4265 264 4267 304
rect 4331 264 4333 304
rect 4337 264 4343 304
rect 4347 264 4349 304
rect 4403 264 4405 304
rect 4409 264 4411 304
rect 4423 264 4425 304
rect 4429 292 4445 304
rect 4429 264 4431 292
rect 4443 264 4445 292
rect 4449 264 4451 304
rect 4503 264 4505 284
rect 4509 264 4511 284
rect 4549 264 4551 304
rect 4555 284 4568 304
rect 4731 284 4741 304
rect 4555 264 4559 284
rect 4571 264 4573 284
rect 4577 264 4583 284
rect 4587 264 4589 284
rect 4601 264 4603 284
rect 4607 264 4611 284
rect 4615 264 4617 284
rect 4655 264 4657 284
rect 4661 264 4665 284
rect 4677 264 4679 284
rect 4683 264 4689 284
rect 4693 264 4695 284
rect 4707 264 4711 284
rect 4715 264 4721 284
rect 4725 264 4727 284
rect 4739 264 4741 284
rect 4745 264 4747 304
rect 66 178 68 236
rect 54 176 68 178
rect 72 176 76 236
rect 80 176 84 236
rect 88 176 90 236
rect 132 196 134 236
rect 138 196 142 236
rect 146 196 148 236
rect 160 216 164 236
rect 168 216 170 236
rect 243 196 245 236
rect 249 196 251 236
rect 263 196 265 236
rect 269 208 271 236
rect 283 208 285 236
rect 269 196 285 208
rect 289 196 291 236
rect 329 196 331 236
rect 335 208 337 236
rect 349 208 351 236
rect 335 196 351 208
rect 355 196 357 236
rect 369 196 371 236
rect 375 196 377 236
rect 466 178 468 236
rect 454 176 468 178
rect 472 176 476 236
rect 480 176 484 236
rect 488 176 490 236
rect 530 176 532 236
rect 536 176 540 236
rect 544 176 548 236
rect 552 178 554 236
rect 632 196 634 236
rect 638 196 642 236
rect 646 196 648 236
rect 660 216 664 236
rect 668 216 670 236
rect 750 216 752 236
rect 756 216 760 236
rect 552 176 566 178
rect 772 196 774 236
rect 778 196 782 236
rect 786 196 788 236
rect 829 216 831 236
rect 835 216 837 236
rect 903 196 905 236
rect 909 196 911 236
rect 923 196 925 236
rect 929 208 931 236
rect 943 208 945 236
rect 929 196 945 208
rect 949 196 951 236
rect 1003 216 1005 236
rect 1009 216 1011 236
rect 1049 196 1051 236
rect 1055 208 1057 236
rect 1069 208 1071 236
rect 1055 196 1071 208
rect 1075 196 1077 236
rect 1089 196 1091 236
rect 1095 196 1097 236
rect 1149 196 1151 236
rect 1155 208 1157 236
rect 1169 208 1171 236
rect 1155 196 1171 208
rect 1175 196 1177 236
rect 1189 196 1191 236
rect 1195 196 1197 236
rect 1250 176 1252 236
rect 1256 176 1260 236
rect 1264 176 1268 236
rect 1272 178 1274 236
rect 1272 176 1286 178
rect 1350 176 1352 236
rect 1356 176 1360 236
rect 1364 176 1368 236
rect 1372 178 1374 236
rect 1470 216 1472 236
rect 1476 216 1480 236
rect 1372 176 1386 178
rect 1492 196 1494 236
rect 1498 196 1502 236
rect 1506 196 1508 236
rect 1550 176 1552 236
rect 1556 176 1560 236
rect 1564 176 1568 236
rect 1572 178 1574 236
rect 1670 216 1672 236
rect 1676 216 1680 236
rect 1572 176 1586 178
rect 1692 196 1694 236
rect 1698 196 1702 236
rect 1706 196 1708 236
rect 1750 176 1752 236
rect 1756 176 1760 236
rect 1764 176 1768 236
rect 1772 178 1774 236
rect 1851 196 1853 236
rect 1857 196 1863 236
rect 1867 196 1869 236
rect 1929 216 1931 236
rect 1935 216 1939 236
rect 1772 176 1786 178
rect 1951 196 1953 236
rect 1957 196 1959 236
rect 2033 196 2035 236
rect 2039 196 2041 236
rect 2053 196 2055 236
rect 2059 196 2065 236
rect 2069 196 2071 236
rect 2109 216 2111 236
rect 2115 216 2119 236
rect 2131 196 2133 236
rect 2137 196 2139 236
rect 2190 176 2192 236
rect 2196 176 2200 236
rect 2204 176 2208 236
rect 2212 178 2214 236
rect 2292 196 2294 236
rect 2298 196 2302 236
rect 2306 196 2308 236
rect 2320 196 2322 236
rect 2326 196 2330 236
rect 2334 196 2336 236
rect 2409 196 2411 236
rect 2415 208 2417 236
rect 2429 208 2431 236
rect 2415 196 2431 208
rect 2435 196 2437 236
rect 2449 196 2451 236
rect 2455 196 2457 236
rect 2530 216 2532 236
rect 2536 216 2540 236
rect 2212 176 2226 178
rect 2552 196 2554 236
rect 2558 196 2562 236
rect 2566 196 2568 236
rect 2609 196 2611 236
rect 2615 208 2617 236
rect 2629 208 2631 236
rect 2615 196 2631 208
rect 2635 196 2637 236
rect 2649 196 2651 236
rect 2655 196 2657 236
rect 2709 216 2711 236
rect 2715 216 2717 236
rect 2770 176 2772 236
rect 2776 176 2780 236
rect 2784 176 2788 236
rect 2792 178 2794 236
rect 2869 216 2871 236
rect 2875 216 2877 236
rect 2792 176 2806 178
rect 2933 196 2935 236
rect 2939 216 2941 236
rect 2953 216 2955 236
rect 2959 216 2965 236
rect 2969 216 2973 236
rect 2985 216 2987 236
rect 2991 216 2997 236
rect 3001 216 3003 236
rect 3015 216 3019 236
rect 3023 216 3025 236
rect 3063 216 3065 236
rect 3069 216 3073 236
rect 3077 216 3079 236
rect 3091 216 3093 236
rect 3097 216 3103 236
rect 3107 216 3109 236
rect 3121 216 3125 236
rect 2939 196 2949 216
rect 3112 196 3125 216
rect 3129 196 3131 236
rect 3169 216 3171 236
rect 3175 216 3177 236
rect 3243 216 3245 236
rect 3249 216 3251 236
rect 3293 196 3295 236
rect 3299 216 3301 236
rect 3313 216 3315 236
rect 3319 216 3325 236
rect 3329 216 3333 236
rect 3345 216 3347 236
rect 3351 216 3357 236
rect 3361 216 3363 236
rect 3375 216 3379 236
rect 3383 216 3385 236
rect 3423 216 3425 236
rect 3429 216 3433 236
rect 3437 216 3439 236
rect 3451 216 3453 236
rect 3457 216 3463 236
rect 3467 216 3469 236
rect 3481 216 3485 236
rect 3299 196 3309 216
rect 3472 196 3485 216
rect 3489 196 3491 236
rect 3543 216 3545 236
rect 3549 216 3551 236
rect 3563 216 3565 236
rect 3569 216 3571 236
rect 3609 196 3611 236
rect 3615 216 3619 236
rect 3631 216 3633 236
rect 3637 216 3643 236
rect 3647 216 3649 236
rect 3661 216 3663 236
rect 3667 216 3671 236
rect 3675 216 3677 236
rect 3715 216 3717 236
rect 3721 216 3725 236
rect 3737 216 3739 236
rect 3743 216 3749 236
rect 3753 216 3755 236
rect 3767 216 3771 236
rect 3775 216 3781 236
rect 3785 216 3787 236
rect 3799 216 3801 236
rect 3615 196 3628 216
rect 3791 196 3801 216
rect 3805 196 3807 236
rect 3849 216 3851 236
rect 3855 216 3857 236
rect 3909 196 3911 236
rect 3915 208 3917 236
rect 3929 208 3931 236
rect 3915 196 3931 208
rect 3935 196 3937 236
rect 3949 196 3951 236
rect 3955 196 3957 236
rect 4009 216 4011 236
rect 4015 216 4017 236
rect 4029 216 4031 236
rect 4035 216 4037 236
rect 4089 216 4091 236
rect 4095 216 4097 236
rect 4109 216 4111 236
rect 4115 216 4117 236
rect 4183 216 4185 236
rect 4189 216 4191 236
rect 4203 216 4205 236
rect 4209 216 4211 236
rect 4249 196 4251 236
rect 4255 208 4257 236
rect 4269 208 4271 236
rect 4255 196 4271 208
rect 4275 196 4277 236
rect 4289 196 4291 236
rect 4295 196 4297 236
rect 4371 196 4373 236
rect 4377 196 4383 236
rect 4387 196 4389 236
rect 4443 216 4445 236
rect 4449 216 4451 236
rect 4489 216 4491 236
rect 4495 216 4497 236
rect 4509 216 4511 236
rect 4515 216 4517 236
rect 4571 196 4573 236
rect 4577 196 4583 236
rect 4587 196 4589 236
rect 4663 216 4665 236
rect 4669 216 4671 236
rect 4711 196 4713 236
rect 4717 196 4723 236
rect 4727 196 4729 236
<< pdiffusion >>
rect 43 4344 45 4424
rect 49 4344 51 4424
rect 63 4344 65 4424
rect 69 4412 85 4424
rect 69 4344 71 4412
rect 83 4344 85 4412
rect 89 4416 103 4424
rect 89 4344 91 4416
rect 417 4416 431 4424
rect 143 4344 145 4384
rect 149 4380 165 4384
rect 149 4344 151 4380
rect 163 4344 165 4380
rect 169 4344 171 4384
rect 183 4344 185 4384
rect 189 4344 191 4384
rect 229 4344 231 4384
rect 235 4344 237 4384
rect 249 4344 251 4384
rect 255 4380 271 4384
rect 255 4344 257 4380
rect 269 4344 271 4380
rect 275 4344 277 4384
rect 343 4344 345 4384
rect 349 4380 365 4384
rect 349 4344 351 4380
rect 363 4344 365 4380
rect 369 4344 371 4384
rect 383 4344 385 4384
rect 389 4344 391 4384
rect 429 4344 431 4416
rect 435 4412 451 4424
rect 435 4344 437 4412
rect 449 4344 451 4412
rect 455 4344 457 4424
rect 469 4344 471 4424
rect 475 4344 477 4424
rect 534 4344 536 4424
rect 540 4344 544 4424
rect 548 4344 550 4424
rect 562 4344 566 4384
rect 570 4344 572 4384
rect 634 4344 636 4424
rect 640 4344 644 4424
rect 648 4344 650 4424
rect 1097 4416 1111 4424
rect 662 4344 666 4384
rect 670 4344 672 4384
rect 743 4344 745 4384
rect 749 4380 765 4384
rect 749 4344 751 4380
rect 763 4344 765 4380
rect 769 4344 771 4384
rect 783 4344 785 4384
rect 789 4344 791 4384
rect 829 4344 831 4384
rect 835 4344 837 4384
rect 849 4344 851 4384
rect 855 4380 871 4384
rect 855 4344 857 4380
rect 869 4344 871 4380
rect 875 4344 877 4384
rect 929 4344 931 4384
rect 935 4344 937 4384
rect 949 4344 951 4384
rect 955 4344 957 4384
rect 1009 4344 1011 4384
rect 1015 4344 1017 4384
rect 1029 4344 1031 4384
rect 1035 4380 1051 4384
rect 1035 4344 1037 4380
rect 1049 4344 1051 4380
rect 1055 4344 1057 4384
rect 1109 4344 1111 4416
rect 1115 4412 1131 4424
rect 1115 4344 1117 4412
rect 1129 4344 1131 4412
rect 1135 4344 1137 4424
rect 1149 4344 1151 4424
rect 1155 4344 1157 4424
rect 1223 4344 1225 4384
rect 1229 4344 1231 4384
rect 1243 4344 1245 4384
rect 1249 4344 1251 4384
rect 1315 4344 1317 4424
rect 1321 4344 1325 4424
rect 1329 4344 1331 4424
rect 1388 4344 1390 4384
rect 1394 4344 1398 4384
rect 1410 4344 1412 4424
rect 1416 4344 1420 4424
rect 1424 4344 1426 4424
rect 1483 4344 1485 4384
rect 1489 4344 1491 4384
rect 1503 4344 1505 4384
rect 1509 4344 1511 4384
rect 1549 4344 1551 4424
rect 1555 4344 1559 4424
rect 1563 4344 1565 4424
rect 1629 4344 1631 4384
rect 1635 4344 1637 4384
rect 1649 4344 1651 4384
rect 1655 4380 1671 4384
rect 1655 4344 1657 4380
rect 1669 4344 1671 4380
rect 1675 4344 1677 4384
rect 1743 4344 1745 4424
rect 1749 4344 1751 4424
rect 1763 4344 1765 4424
rect 1769 4412 1785 4424
rect 1769 4344 1771 4412
rect 1783 4344 1785 4412
rect 1789 4416 1803 4424
rect 1789 4344 1791 4416
rect 1937 4416 1951 4424
rect 1829 4344 1831 4384
rect 1835 4344 1837 4384
rect 1903 4344 1905 4384
rect 1909 4344 1911 4384
rect 1949 4344 1951 4416
rect 1955 4412 1971 4424
rect 1955 4344 1957 4412
rect 1969 4344 1971 4412
rect 1975 4344 1977 4424
rect 1989 4344 1991 4424
rect 1995 4344 1997 4424
rect 2049 4344 2051 4424
rect 2055 4344 2059 4424
rect 2063 4344 2065 4424
rect 2129 4344 2131 4384
rect 2135 4344 2137 4384
rect 2194 4344 2196 4424
rect 2200 4344 2204 4424
rect 2208 4344 2210 4424
rect 2222 4344 2226 4384
rect 2230 4344 2232 4384
rect 2313 4344 2315 4424
rect 2319 4344 2325 4424
rect 2329 4344 2331 4424
rect 2353 4344 2355 4424
rect 2359 4344 2365 4424
rect 2369 4344 2371 4424
rect 2409 4344 2411 4424
rect 2415 4344 2421 4424
rect 2425 4423 2441 4424
rect 2425 4344 2427 4423
rect 2439 4344 2441 4423
rect 2445 4423 2459 4424
rect 2445 4344 2447 4423
rect 2497 4416 2511 4424
rect 2509 4344 2511 4416
rect 2515 4412 2531 4424
rect 2515 4344 2517 4412
rect 2529 4344 2531 4412
rect 2535 4344 2537 4424
rect 2549 4344 2551 4424
rect 2555 4344 2557 4424
rect 2623 4344 2625 4424
rect 2629 4356 2631 4424
rect 2643 4356 2645 4424
rect 2629 4344 2645 4356
rect 2649 4422 2665 4424
rect 2649 4344 2651 4422
rect 2663 4344 2665 4422
rect 2669 4410 2685 4424
rect 2669 4344 2671 4410
rect 2683 4344 2685 4410
rect 2689 4422 2703 4424
rect 2689 4344 2691 4422
rect 2733 4344 2735 4424
rect 2739 4384 2748 4424
rect 2739 4344 2741 4384
rect 2753 4344 2755 4384
rect 2759 4344 2769 4384
rect 2773 4344 2775 4384
rect 2787 4344 2789 4384
rect 2793 4344 2801 4384
rect 2805 4344 2807 4384
rect 2819 4344 2821 4384
rect 2825 4344 2827 4384
rect 2865 4344 2867 4384
rect 2871 4344 2875 4384
rect 2879 4364 2890 4384
rect 2916 4364 2925 4424
rect 2879 4344 2881 4364
rect 2893 4344 2895 4364
rect 2899 4344 2903 4364
rect 2907 4344 2911 4364
rect 2923 4344 2925 4364
rect 2929 4344 2931 4424
rect 2983 4344 2985 4384
rect 2989 4344 2991 4384
rect 3048 4344 3050 4384
rect 3054 4344 3058 4384
rect 3070 4344 3072 4424
rect 3076 4344 3080 4424
rect 3084 4344 3086 4424
rect 3155 4344 3157 4424
rect 3161 4344 3165 4424
rect 3169 4344 3171 4424
rect 3228 4344 3230 4384
rect 3234 4344 3238 4384
rect 3250 4344 3252 4424
rect 3256 4344 3260 4424
rect 3264 4344 3266 4424
rect 3335 4344 3337 4424
rect 3341 4344 3345 4424
rect 3349 4344 3351 4424
rect 3403 4344 3405 4384
rect 3409 4344 3411 4384
rect 3449 4344 3451 4424
rect 3455 4364 3464 4424
rect 3632 4384 3641 4424
rect 3490 4364 3501 4384
rect 3455 4344 3457 4364
rect 3469 4344 3473 4364
rect 3477 4344 3481 4364
rect 3485 4344 3487 4364
rect 3499 4344 3501 4364
rect 3505 4344 3509 4384
rect 3513 4344 3515 4384
rect 3553 4344 3555 4384
rect 3559 4344 3561 4384
rect 3573 4344 3575 4384
rect 3579 4344 3587 4384
rect 3591 4344 3593 4384
rect 3605 4344 3607 4384
rect 3611 4344 3621 4384
rect 3625 4344 3627 4384
rect 3639 4344 3641 4384
rect 3645 4344 3647 4424
rect 3694 4344 3696 4424
rect 3700 4344 3704 4424
rect 3708 4344 3710 4424
rect 3722 4344 3726 4384
rect 3730 4344 3732 4384
rect 3789 4344 3791 4384
rect 3795 4344 3797 4384
rect 3809 4344 3811 4384
rect 3815 4344 3817 4384
rect 3883 4344 3885 4424
rect 3889 4344 3891 4424
rect 3903 4344 3905 4424
rect 3909 4344 3911 4424
rect 3923 4344 3925 4424
rect 3929 4344 3931 4424
rect 3943 4344 3945 4424
rect 3949 4344 3951 4424
rect 3963 4344 3965 4424
rect 3969 4344 3971 4424
rect 3983 4344 3985 4424
rect 3989 4344 3991 4424
rect 4003 4344 4005 4424
rect 4009 4344 4011 4424
rect 4023 4344 4025 4424
rect 4029 4344 4031 4424
rect 4081 4344 4083 4424
rect 4087 4344 4089 4424
rect 4101 4344 4105 4384
rect 4109 4344 4111 4384
rect 4149 4344 4151 4384
rect 4155 4344 4157 4384
rect 4169 4344 4171 4384
rect 4175 4344 4177 4384
rect 4229 4344 4231 4384
rect 4235 4344 4237 4384
rect 4294 4344 4296 4424
rect 4300 4344 4304 4424
rect 4308 4344 4310 4424
rect 4322 4344 4326 4384
rect 4330 4344 4332 4384
rect 4389 4344 4391 4424
rect 4395 4364 4404 4424
rect 4572 4384 4581 4424
rect 4430 4364 4441 4384
rect 4395 4344 4397 4364
rect 4409 4344 4413 4364
rect 4417 4344 4421 4364
rect 4425 4344 4427 4364
rect 4439 4344 4441 4364
rect 4445 4344 4449 4384
rect 4453 4344 4455 4384
rect 4493 4344 4495 4384
rect 4499 4344 4501 4384
rect 4513 4344 4515 4384
rect 4519 4344 4527 4384
rect 4531 4344 4533 4384
rect 4545 4344 4547 4384
rect 4551 4344 4561 4384
rect 4565 4344 4567 4384
rect 4579 4344 4581 4384
rect 4585 4344 4587 4424
rect 4629 4344 4631 4384
rect 4635 4344 4639 4384
rect 4651 4344 4653 4424
rect 4657 4344 4659 4424
rect 4709 4344 4711 4384
rect 4715 4344 4717 4384
rect 4729 4344 4731 4384
rect 4735 4344 4737 4384
rect 43 4276 45 4316
rect 49 4276 51 4316
rect 63 4276 65 4316
rect 69 4276 71 4316
rect 109 4244 111 4316
rect 97 4236 111 4244
rect 115 4248 117 4316
rect 129 4248 131 4316
rect 115 4236 131 4248
rect 135 4236 137 4316
rect 149 4236 151 4316
rect 155 4236 157 4316
rect 223 4276 225 4316
rect 229 4276 231 4316
rect 243 4276 245 4316
rect 249 4276 251 4316
rect 315 4236 317 4316
rect 321 4236 325 4316
rect 329 4236 331 4316
rect 388 4276 390 4316
rect 394 4276 398 4316
rect 410 4236 412 4316
rect 416 4236 420 4316
rect 424 4236 426 4316
rect 474 4236 476 4316
rect 480 4236 484 4316
rect 488 4236 490 4316
rect 502 4276 506 4316
rect 510 4276 512 4316
rect 583 4276 585 4316
rect 589 4276 591 4316
rect 643 4236 645 4316
rect 649 4236 651 4316
rect 663 4236 665 4316
rect 669 4248 671 4316
rect 683 4248 685 4316
rect 669 4236 685 4248
rect 689 4244 691 4316
rect 743 4276 745 4316
rect 749 4276 751 4316
rect 789 4276 791 4316
rect 795 4276 797 4316
rect 809 4276 811 4316
rect 815 4280 817 4316
rect 829 4280 831 4316
rect 815 4276 831 4280
rect 835 4276 837 4316
rect 689 4236 703 4244
rect 903 4236 905 4316
rect 909 4304 925 4316
rect 909 4236 911 4304
rect 923 4236 925 4304
rect 929 4238 931 4316
rect 943 4238 945 4316
rect 929 4236 945 4238
rect 949 4250 951 4316
rect 963 4250 965 4316
rect 949 4236 965 4250
rect 969 4238 971 4316
rect 1023 4276 1025 4316
rect 1029 4280 1031 4316
rect 1043 4280 1045 4316
rect 1029 4276 1045 4280
rect 1049 4276 1051 4316
rect 1063 4276 1065 4316
rect 1069 4276 1071 4316
rect 1109 4276 1111 4316
rect 1115 4276 1117 4316
rect 1129 4276 1131 4316
rect 1135 4280 1137 4316
rect 1149 4280 1151 4316
rect 1135 4276 1151 4280
rect 1155 4276 1157 4316
rect 1223 4276 1225 4316
rect 1229 4276 1231 4316
rect 1243 4276 1245 4316
rect 1249 4276 1251 4316
rect 1303 4276 1305 4316
rect 1309 4280 1311 4316
rect 1323 4280 1325 4316
rect 1309 4276 1325 4280
rect 1329 4276 1331 4316
rect 1343 4276 1345 4316
rect 1349 4276 1351 4316
rect 1403 4276 1405 4316
rect 1409 4276 1411 4316
rect 1423 4276 1425 4316
rect 1429 4276 1431 4316
rect 1469 4276 1471 4316
rect 1475 4276 1477 4316
rect 1489 4276 1491 4316
rect 1495 4280 1497 4316
rect 1509 4280 1511 4316
rect 1495 4276 1511 4280
rect 1515 4276 1517 4316
rect 969 4236 983 4238
rect 1595 4236 1597 4316
rect 1601 4236 1605 4316
rect 1609 4236 1611 4316
rect 1675 4236 1677 4316
rect 1681 4236 1685 4316
rect 1689 4236 1691 4316
rect 1734 4236 1736 4316
rect 1740 4236 1744 4316
rect 1748 4236 1750 4316
rect 1762 4276 1766 4316
rect 1770 4276 1772 4316
rect 1843 4276 1845 4316
rect 1849 4276 1851 4316
rect 1863 4276 1865 4316
rect 1869 4276 1871 4316
rect 1909 4276 1911 4316
rect 1915 4276 1917 4316
rect 1969 4276 1971 4316
rect 1975 4276 1977 4316
rect 1989 4276 1991 4316
rect 1995 4280 1997 4316
rect 2009 4280 2011 4316
rect 1995 4276 2011 4280
rect 2015 4276 2017 4316
rect 2069 4276 2071 4316
rect 2075 4276 2077 4316
rect 2089 4276 2091 4316
rect 2095 4280 2097 4316
rect 2109 4280 2111 4316
rect 2095 4276 2111 4280
rect 2115 4276 2117 4316
rect 2173 4236 2175 4316
rect 2179 4276 2181 4316
rect 2193 4276 2195 4316
rect 2199 4276 2209 4316
rect 2213 4276 2215 4316
rect 2227 4276 2229 4316
rect 2233 4276 2241 4316
rect 2245 4276 2247 4316
rect 2259 4276 2261 4316
rect 2265 4276 2267 4316
rect 2305 4276 2307 4316
rect 2311 4276 2315 4316
rect 2319 4296 2321 4316
rect 2333 4296 2335 4316
rect 2339 4296 2343 4316
rect 2347 4296 2351 4316
rect 2363 4296 2365 4316
rect 2319 4276 2330 4296
rect 2179 4236 2188 4276
rect 2356 4236 2365 4296
rect 2369 4236 2371 4316
rect 2409 4276 2411 4316
rect 2415 4276 2419 4316
rect 2431 4236 2433 4316
rect 2437 4236 2439 4316
rect 2503 4276 2505 4316
rect 2509 4276 2511 4316
rect 2575 4236 2577 4316
rect 2581 4236 2585 4316
rect 2589 4236 2591 4316
rect 2629 4236 2631 4316
rect 2635 4296 2637 4316
rect 2649 4296 2653 4316
rect 2657 4296 2661 4316
rect 2665 4296 2667 4316
rect 2679 4296 2681 4316
rect 2635 4236 2644 4296
rect 2670 4276 2681 4296
rect 2685 4276 2689 4316
rect 2693 4276 2695 4316
rect 2733 4276 2735 4316
rect 2739 4276 2741 4316
rect 2753 4276 2755 4316
rect 2759 4276 2767 4316
rect 2771 4276 2773 4316
rect 2785 4276 2787 4316
rect 2791 4276 2801 4316
rect 2805 4276 2807 4316
rect 2819 4276 2821 4316
rect 2812 4236 2821 4276
rect 2825 4236 2827 4316
rect 2869 4276 2871 4316
rect 2875 4276 2877 4316
rect 2955 4236 2957 4316
rect 2961 4236 2965 4316
rect 2969 4236 2971 4316
rect 3014 4236 3016 4316
rect 3020 4236 3024 4316
rect 3028 4236 3030 4316
rect 3042 4276 3046 4316
rect 3050 4276 3052 4316
rect 3109 4276 3111 4316
rect 3115 4276 3117 4316
rect 3129 4276 3131 4316
rect 3135 4276 3137 4316
rect 3203 4276 3205 4316
rect 3209 4276 3211 4316
rect 3223 4276 3225 4316
rect 3229 4276 3231 4316
rect 3283 4276 3285 4316
rect 3289 4276 3291 4316
rect 3303 4276 3305 4316
rect 3309 4276 3311 4316
rect 3349 4236 3351 4316
rect 3355 4236 3359 4316
rect 3363 4236 3365 4316
rect 3433 4236 3435 4316
rect 3439 4276 3441 4316
rect 3453 4276 3455 4316
rect 3459 4276 3469 4316
rect 3473 4276 3475 4316
rect 3487 4276 3489 4316
rect 3493 4276 3501 4316
rect 3505 4276 3507 4316
rect 3519 4276 3521 4316
rect 3525 4276 3527 4316
rect 3565 4276 3567 4316
rect 3571 4276 3575 4316
rect 3579 4296 3581 4316
rect 3593 4296 3595 4316
rect 3599 4296 3603 4316
rect 3607 4296 3611 4316
rect 3623 4296 3625 4316
rect 3579 4276 3590 4296
rect 3439 4236 3448 4276
rect 3616 4236 3625 4296
rect 3629 4236 3631 4316
rect 3683 4276 3685 4316
rect 3689 4276 3691 4316
rect 3703 4276 3705 4316
rect 3709 4276 3711 4316
rect 3749 4236 3751 4316
rect 3755 4236 3759 4316
rect 3763 4236 3765 4316
rect 3829 4236 3831 4316
rect 3835 4296 3837 4316
rect 3849 4296 3853 4316
rect 3857 4296 3861 4316
rect 3865 4296 3867 4316
rect 3879 4296 3881 4316
rect 3835 4236 3844 4296
rect 3870 4276 3881 4296
rect 3885 4276 3889 4316
rect 3893 4276 3895 4316
rect 3933 4276 3935 4316
rect 3939 4276 3941 4316
rect 3953 4276 3955 4316
rect 3959 4276 3967 4316
rect 3971 4276 3973 4316
rect 3985 4276 3987 4316
rect 3991 4276 4001 4316
rect 4005 4276 4007 4316
rect 4019 4276 4021 4316
rect 4012 4236 4021 4276
rect 4025 4236 4027 4316
rect 4069 4236 4071 4316
rect 4075 4236 4079 4316
rect 4083 4236 4085 4316
rect 4163 4236 4165 4316
rect 4169 4236 4171 4316
rect 4183 4236 4185 4316
rect 4189 4248 4191 4316
rect 4203 4248 4205 4316
rect 4189 4236 4205 4248
rect 4209 4244 4211 4316
rect 4249 4276 4251 4316
rect 4255 4276 4259 4316
rect 4209 4236 4223 4244
rect 4271 4236 4273 4316
rect 4277 4236 4279 4316
rect 4355 4236 4357 4316
rect 4361 4236 4365 4316
rect 4369 4236 4371 4316
rect 4423 4236 4425 4316
rect 4429 4236 4431 4316
rect 4443 4236 4445 4316
rect 4449 4248 4451 4316
rect 4463 4248 4465 4316
rect 4449 4236 4465 4248
rect 4469 4244 4471 4316
rect 4469 4236 4483 4244
rect 4509 4236 4511 4316
rect 4515 4296 4517 4316
rect 4529 4296 4533 4316
rect 4537 4296 4541 4316
rect 4545 4296 4547 4316
rect 4559 4296 4561 4316
rect 4515 4236 4524 4296
rect 4550 4276 4561 4296
rect 4565 4276 4569 4316
rect 4573 4276 4575 4316
rect 4613 4276 4615 4316
rect 4619 4276 4621 4316
rect 4633 4276 4635 4316
rect 4639 4276 4647 4316
rect 4651 4276 4653 4316
rect 4665 4276 4667 4316
rect 4671 4276 4681 4316
rect 4685 4276 4687 4316
rect 4699 4276 4701 4316
rect 4692 4236 4701 4276
rect 4705 4236 4707 4316
rect 43 3864 45 3904
rect 49 3864 51 3904
rect 63 3864 65 3904
rect 69 3864 71 3904
rect 109 3864 111 3904
rect 115 3864 117 3904
rect 129 3864 131 3904
rect 135 3864 137 3904
rect 203 3864 205 3904
rect 209 3864 211 3904
rect 223 3864 225 3904
rect 229 3864 231 3904
rect 288 3864 290 3904
rect 294 3864 298 3904
rect 310 3864 312 3944
rect 316 3864 320 3944
rect 324 3864 326 3944
rect 357 3936 371 3944
rect 369 3864 371 3936
rect 375 3932 391 3944
rect 375 3864 377 3932
rect 389 3864 391 3932
rect 395 3864 397 3944
rect 409 3864 411 3944
rect 415 3864 417 3944
rect 495 3864 497 3944
rect 501 3864 505 3944
rect 509 3864 511 3944
rect 549 3864 551 3904
rect 555 3864 557 3904
rect 569 3864 571 3904
rect 575 3864 577 3904
rect 634 3864 636 3944
rect 640 3864 644 3944
rect 648 3864 650 3944
rect 662 3864 666 3904
rect 670 3864 672 3904
rect 743 3864 745 3904
rect 749 3900 765 3904
rect 749 3864 751 3900
rect 763 3864 765 3900
rect 769 3864 771 3904
rect 783 3864 785 3904
rect 789 3864 791 3904
rect 829 3864 831 3904
rect 835 3864 837 3904
rect 849 3864 851 3904
rect 855 3900 871 3904
rect 855 3864 857 3900
rect 869 3864 871 3900
rect 875 3864 877 3904
rect 948 3864 950 3904
rect 954 3864 958 3904
rect 970 3864 972 3944
rect 976 3864 980 3944
rect 984 3864 986 3944
rect 1034 3864 1036 3944
rect 1040 3864 1044 3944
rect 1048 3864 1050 3944
rect 1062 3864 1066 3904
rect 1070 3864 1072 3904
rect 1143 3864 1145 3904
rect 1149 3864 1151 3904
rect 1203 3864 1205 3904
rect 1209 3900 1225 3904
rect 1209 3864 1211 3900
rect 1223 3864 1225 3900
rect 1229 3864 1231 3904
rect 1243 3864 1245 3904
rect 1249 3864 1251 3904
rect 1289 3864 1291 3904
rect 1295 3864 1297 3904
rect 1349 3864 1351 3904
rect 1355 3864 1357 3904
rect 1369 3864 1371 3904
rect 1375 3900 1391 3904
rect 1375 3864 1377 3900
rect 1389 3864 1391 3900
rect 1395 3864 1397 3904
rect 1449 3864 1451 3904
rect 1455 3864 1457 3904
rect 1469 3864 1471 3904
rect 1475 3900 1491 3904
rect 1475 3864 1477 3900
rect 1489 3864 1491 3900
rect 1495 3864 1497 3904
rect 1549 3864 1551 3904
rect 1555 3864 1557 3904
rect 1569 3864 1571 3904
rect 1575 3864 1577 3904
rect 1655 3864 1657 3944
rect 1661 3864 1665 3944
rect 1669 3864 1671 3944
rect 1719 3864 1721 3944
rect 1725 3864 1727 3944
rect 1739 3864 1743 3904
rect 1747 3864 1751 3904
rect 1763 3864 1765 3904
rect 1769 3864 1771 3904
rect 1828 3864 1830 3904
rect 1834 3864 1838 3904
rect 1850 3864 1852 3944
rect 1856 3864 1860 3944
rect 1864 3864 1866 3944
rect 1909 3864 1911 3944
rect 1915 3864 1919 3944
rect 1923 3864 1925 3944
rect 2003 3864 2005 3904
rect 2009 3864 2011 3904
rect 2054 3864 2056 3944
rect 2060 3864 2064 3944
rect 2068 3864 2070 3944
rect 2082 3864 2086 3904
rect 2090 3864 2092 3904
rect 2149 3864 2151 3904
rect 2155 3864 2157 3904
rect 2209 3864 2211 3904
rect 2215 3864 2217 3904
rect 2229 3864 2231 3904
rect 2235 3864 2237 3904
rect 2289 3864 2291 3904
rect 2295 3864 2297 3904
rect 2309 3864 2311 3904
rect 2315 3900 2331 3904
rect 2315 3864 2317 3900
rect 2329 3864 2331 3900
rect 2335 3864 2337 3904
rect 2389 3864 2391 3904
rect 2395 3864 2399 3904
rect 2411 3864 2413 3944
rect 2417 3864 2419 3944
rect 2469 3864 2471 3944
rect 2475 3864 2477 3944
rect 2489 3864 2491 3944
rect 2495 3864 2497 3944
rect 2509 3864 2511 3944
rect 2515 3864 2517 3944
rect 2529 3864 2531 3944
rect 2535 3864 2537 3944
rect 2549 3864 2551 3944
rect 2555 3864 2557 3944
rect 2569 3864 2571 3944
rect 2575 3864 2577 3944
rect 2589 3864 2591 3944
rect 2595 3864 2597 3944
rect 2609 3864 2611 3944
rect 2615 3864 2617 3944
rect 2673 3864 2675 3944
rect 2679 3904 2688 3944
rect 2679 3864 2681 3904
rect 2693 3864 2695 3904
rect 2699 3864 2709 3904
rect 2713 3864 2715 3904
rect 2727 3864 2729 3904
rect 2733 3864 2741 3904
rect 2745 3864 2747 3904
rect 2759 3864 2761 3904
rect 2765 3864 2767 3904
rect 2805 3864 2807 3904
rect 2811 3864 2815 3904
rect 2819 3884 2830 3904
rect 2856 3884 2865 3944
rect 2819 3864 2821 3884
rect 2833 3864 2835 3884
rect 2839 3864 2843 3884
rect 2847 3864 2851 3884
rect 2863 3864 2865 3884
rect 2869 3864 2871 3944
rect 2909 3864 2911 3904
rect 2915 3864 2917 3904
rect 2974 3864 2976 3944
rect 2980 3864 2984 3944
rect 2988 3864 2990 3944
rect 3002 3864 3006 3904
rect 3010 3864 3012 3904
rect 3069 3864 3071 3944
rect 3075 3864 3079 3944
rect 3083 3864 3085 3944
rect 3149 3864 3151 3904
rect 3155 3864 3157 3904
rect 3169 3864 3171 3904
rect 3175 3864 3177 3904
rect 3243 3864 3245 3944
rect 3249 3864 3251 3944
rect 3263 3864 3265 3944
rect 3269 3932 3285 3944
rect 3269 3864 3271 3932
rect 3283 3864 3285 3932
rect 3289 3936 3303 3944
rect 3289 3864 3291 3936
rect 3329 3864 3331 3904
rect 3335 3864 3337 3904
rect 3349 3864 3353 3904
rect 3357 3864 3361 3904
rect 3373 3864 3375 3944
rect 3379 3864 3381 3944
rect 3455 3864 3457 3944
rect 3461 3864 3465 3944
rect 3469 3864 3471 3944
rect 3523 3864 3525 3904
rect 3529 3864 3531 3904
rect 3569 3864 3571 3944
rect 3575 3884 3584 3944
rect 3752 3904 3761 3944
rect 3610 3884 3621 3904
rect 3575 3864 3577 3884
rect 3589 3864 3593 3884
rect 3597 3864 3601 3884
rect 3605 3864 3607 3884
rect 3619 3864 3621 3884
rect 3625 3864 3629 3904
rect 3633 3864 3635 3904
rect 3673 3864 3675 3904
rect 3679 3864 3681 3904
rect 3693 3864 3695 3904
rect 3699 3864 3707 3904
rect 3711 3864 3713 3904
rect 3725 3864 3727 3904
rect 3731 3864 3741 3904
rect 3745 3864 3747 3904
rect 3759 3864 3761 3904
rect 3765 3864 3767 3944
rect 3823 3864 3825 3944
rect 3829 3864 3831 3944
rect 3843 3864 3845 3944
rect 3849 3932 3865 3944
rect 3849 3864 3851 3932
rect 3863 3864 3865 3932
rect 3869 3936 3883 3944
rect 3869 3864 3871 3936
rect 3909 3864 3911 3944
rect 3915 3864 3919 3944
rect 3923 3864 3925 3944
rect 4015 3864 4017 3944
rect 4021 3864 4025 3944
rect 4029 3864 4031 3944
rect 4069 3864 4071 3904
rect 4075 3864 4077 3904
rect 4089 3864 4093 3904
rect 4097 3864 4101 3904
rect 4113 3864 4115 3944
rect 4119 3864 4121 3944
rect 4174 3864 4176 3944
rect 4180 3864 4184 3944
rect 4188 3864 4190 3944
rect 4202 3864 4206 3904
rect 4210 3864 4212 3904
rect 4288 3864 4290 3904
rect 4294 3864 4298 3904
rect 4310 3864 4312 3944
rect 4316 3864 4320 3944
rect 4324 3864 4326 3944
rect 4383 3864 4385 3904
rect 4389 3864 4391 3904
rect 4429 3864 4431 3944
rect 4435 3884 4444 3944
rect 4612 3904 4621 3944
rect 4470 3884 4481 3904
rect 4435 3864 4437 3884
rect 4449 3864 4453 3884
rect 4457 3864 4461 3884
rect 4465 3864 4467 3884
rect 4479 3864 4481 3884
rect 4485 3864 4489 3904
rect 4493 3864 4495 3904
rect 4533 3864 4535 3904
rect 4539 3864 4541 3904
rect 4553 3864 4555 3904
rect 4559 3864 4567 3904
rect 4571 3864 4573 3904
rect 4585 3864 4587 3904
rect 4591 3864 4601 3904
rect 4605 3864 4607 3904
rect 4619 3864 4621 3904
rect 4625 3864 4627 3944
rect 4669 3864 4671 3904
rect 4675 3864 4677 3904
rect 55 3756 57 3836
rect 61 3756 65 3836
rect 69 3756 71 3836
rect 114 3756 116 3836
rect 120 3756 124 3836
rect 128 3756 130 3836
rect 142 3796 146 3836
rect 150 3796 152 3836
rect 223 3796 225 3836
rect 229 3796 231 3836
rect 283 3756 285 3836
rect 289 3756 291 3836
rect 303 3756 305 3836
rect 309 3768 311 3836
rect 323 3768 325 3836
rect 309 3756 325 3768
rect 329 3764 331 3836
rect 329 3756 343 3764
rect 379 3756 381 3836
rect 385 3756 387 3836
rect 399 3796 403 3836
rect 407 3796 411 3836
rect 423 3796 425 3836
rect 429 3796 431 3836
rect 483 3796 485 3836
rect 489 3796 491 3836
rect 503 3796 505 3836
rect 509 3796 511 3836
rect 563 3796 565 3836
rect 569 3796 571 3836
rect 583 3796 585 3836
rect 589 3796 591 3836
rect 629 3796 631 3836
rect 635 3796 637 3836
rect 694 3756 696 3836
rect 700 3756 704 3836
rect 708 3756 710 3836
rect 722 3796 726 3836
rect 730 3796 732 3836
rect 789 3796 791 3836
rect 795 3796 797 3836
rect 809 3796 811 3836
rect 815 3796 817 3836
rect 883 3796 885 3836
rect 889 3800 891 3836
rect 903 3800 905 3836
rect 889 3796 905 3800
rect 909 3796 911 3836
rect 923 3796 925 3836
rect 929 3796 931 3836
rect 969 3764 971 3836
rect 957 3756 971 3764
rect 975 3768 977 3836
rect 989 3768 991 3836
rect 975 3756 991 3768
rect 995 3756 997 3836
rect 1009 3756 1011 3836
rect 1015 3756 1017 3836
rect 1069 3796 1071 3836
rect 1075 3796 1077 3836
rect 1089 3796 1091 3836
rect 1095 3800 1097 3836
rect 1109 3800 1111 3836
rect 1095 3796 1111 3800
rect 1115 3796 1117 3836
rect 1169 3764 1171 3836
rect 1157 3756 1171 3764
rect 1175 3768 1177 3836
rect 1189 3768 1191 3836
rect 1175 3756 1191 3768
rect 1195 3756 1197 3836
rect 1209 3756 1211 3836
rect 1215 3756 1217 3836
rect 1269 3796 1271 3836
rect 1275 3796 1277 3836
rect 1343 3796 1345 3836
rect 1349 3800 1351 3836
rect 1363 3800 1365 3836
rect 1349 3796 1365 3800
rect 1369 3796 1371 3836
rect 1383 3796 1385 3836
rect 1389 3796 1391 3836
rect 1443 3796 1445 3836
rect 1449 3796 1451 3836
rect 1508 3796 1510 3836
rect 1514 3796 1518 3836
rect 1530 3756 1532 3836
rect 1536 3756 1540 3836
rect 1544 3756 1546 3836
rect 1603 3796 1605 3836
rect 1609 3796 1611 3836
rect 1649 3764 1651 3836
rect 1637 3756 1651 3764
rect 1655 3768 1657 3836
rect 1669 3768 1671 3836
rect 1655 3756 1671 3768
rect 1675 3756 1677 3836
rect 1689 3756 1691 3836
rect 1695 3756 1697 3836
rect 1749 3756 1751 3836
rect 1755 3756 1759 3836
rect 1763 3756 1765 3836
rect 1843 3756 1845 3836
rect 1849 3756 1851 3836
rect 1863 3756 1865 3836
rect 1869 3768 1871 3836
rect 1883 3768 1885 3836
rect 1869 3756 1885 3768
rect 1889 3764 1891 3836
rect 1943 3796 1945 3836
rect 1949 3796 1951 3836
rect 1963 3796 1965 3836
rect 1969 3796 1971 3836
rect 1889 3756 1903 3764
rect 2009 3756 2011 3836
rect 2015 3756 2021 3836
rect 2025 3757 2027 3836
rect 2039 3757 2041 3836
rect 2025 3756 2041 3757
rect 2045 3757 2047 3836
rect 2109 3796 2111 3836
rect 2115 3796 2119 3836
rect 2045 3756 2059 3757
rect 2131 3756 2133 3836
rect 2137 3756 2139 3836
rect 2203 3756 2205 3836
rect 2209 3756 2211 3836
rect 2223 3756 2225 3836
rect 2229 3756 2231 3836
rect 2243 3756 2245 3836
rect 2249 3756 2251 3836
rect 2263 3756 2265 3836
rect 2269 3756 2271 3836
rect 2283 3756 2285 3836
rect 2289 3756 2291 3836
rect 2303 3756 2305 3836
rect 2309 3756 2311 3836
rect 2323 3756 2325 3836
rect 2329 3756 2331 3836
rect 2343 3756 2345 3836
rect 2349 3756 2351 3836
rect 2393 3756 2395 3836
rect 2399 3796 2401 3836
rect 2413 3796 2415 3836
rect 2419 3796 2429 3836
rect 2433 3796 2435 3836
rect 2447 3796 2449 3836
rect 2453 3796 2461 3836
rect 2465 3796 2467 3836
rect 2479 3796 2481 3836
rect 2485 3796 2487 3836
rect 2525 3796 2527 3836
rect 2531 3796 2535 3836
rect 2539 3816 2541 3836
rect 2553 3816 2555 3836
rect 2559 3816 2563 3836
rect 2567 3816 2571 3836
rect 2583 3816 2585 3836
rect 2539 3796 2550 3816
rect 2399 3756 2408 3796
rect 2576 3756 2585 3816
rect 2589 3756 2591 3836
rect 2648 3796 2650 3836
rect 2654 3796 2658 3836
rect 2670 3756 2672 3836
rect 2676 3756 2680 3836
rect 2684 3756 2686 3836
rect 2743 3796 2745 3836
rect 2749 3796 2751 3836
rect 2815 3756 2817 3836
rect 2821 3756 2825 3836
rect 2829 3756 2831 3836
rect 2895 3756 2897 3836
rect 2901 3756 2905 3836
rect 2909 3756 2911 3836
rect 2975 3756 2977 3836
rect 2981 3756 2985 3836
rect 2989 3756 2991 3836
rect 3029 3796 3031 3836
rect 3035 3796 3037 3836
rect 3103 3796 3105 3836
rect 3109 3796 3111 3836
rect 3154 3756 3156 3836
rect 3160 3756 3164 3836
rect 3168 3756 3170 3836
rect 3182 3796 3186 3836
rect 3190 3796 3192 3836
rect 3263 3756 3265 3836
rect 3269 3756 3271 3836
rect 3283 3756 3285 3836
rect 3289 3768 3291 3836
rect 3303 3768 3305 3836
rect 3289 3756 3305 3768
rect 3309 3764 3311 3836
rect 3309 3756 3323 3764
rect 3349 3764 3351 3836
rect 3337 3756 3351 3764
rect 3355 3768 3357 3836
rect 3369 3768 3371 3836
rect 3355 3756 3371 3768
rect 3375 3756 3377 3836
rect 3389 3756 3391 3836
rect 3395 3756 3397 3836
rect 3449 3796 3451 3836
rect 3455 3796 3457 3836
rect 3509 3796 3511 3836
rect 3515 3796 3517 3836
rect 3529 3796 3533 3836
rect 3537 3796 3541 3836
rect 3553 3756 3555 3836
rect 3559 3756 3561 3836
rect 3614 3756 3616 3836
rect 3620 3756 3624 3836
rect 3628 3756 3630 3836
rect 3642 3796 3646 3836
rect 3650 3796 3652 3836
rect 3714 3756 3716 3836
rect 3720 3756 3724 3836
rect 3728 3756 3730 3836
rect 3742 3796 3746 3836
rect 3750 3796 3752 3836
rect 3813 3756 3815 3836
rect 3819 3796 3821 3836
rect 3833 3796 3835 3836
rect 3839 3796 3849 3836
rect 3853 3796 3855 3836
rect 3867 3796 3869 3836
rect 3873 3796 3881 3836
rect 3885 3796 3887 3836
rect 3899 3796 3901 3836
rect 3905 3796 3907 3836
rect 3945 3796 3947 3836
rect 3951 3796 3955 3836
rect 3959 3816 3961 3836
rect 3973 3816 3975 3836
rect 3979 3816 3983 3836
rect 3987 3816 3991 3836
rect 4003 3816 4005 3836
rect 3959 3796 3970 3816
rect 3819 3756 3828 3796
rect 3996 3756 4005 3816
rect 4009 3756 4011 3836
rect 4049 3796 4051 3836
rect 4055 3796 4059 3836
rect 4071 3756 4073 3836
rect 4077 3756 4079 3836
rect 4155 3756 4157 3836
rect 4161 3756 4165 3836
rect 4169 3756 4171 3836
rect 4209 3764 4211 3836
rect 4197 3756 4211 3764
rect 4215 3768 4217 3836
rect 4229 3768 4231 3836
rect 4215 3756 4231 3768
rect 4235 3756 4237 3836
rect 4249 3756 4251 3836
rect 4255 3756 4257 3836
rect 4309 3756 4311 3836
rect 4315 3816 4317 3836
rect 4329 3816 4333 3836
rect 4337 3816 4341 3836
rect 4345 3816 4347 3836
rect 4359 3816 4361 3836
rect 4315 3756 4324 3816
rect 4350 3796 4361 3816
rect 4365 3796 4369 3836
rect 4373 3796 4375 3836
rect 4413 3796 4415 3836
rect 4419 3796 4421 3836
rect 4433 3796 4435 3836
rect 4439 3796 4447 3836
rect 4451 3796 4453 3836
rect 4465 3796 4467 3836
rect 4471 3796 4481 3836
rect 4485 3796 4487 3836
rect 4499 3796 4501 3836
rect 4492 3756 4501 3796
rect 4505 3756 4507 3836
rect 4549 3796 4551 3836
rect 4555 3796 4559 3836
rect 4571 3756 4573 3836
rect 4577 3756 4579 3836
rect 4643 3796 4645 3836
rect 4649 3796 4651 3836
rect 4689 3796 4691 3836
rect 4695 3796 4697 3836
rect 43 3384 45 3424
rect 49 3384 51 3424
rect 63 3384 65 3424
rect 69 3384 71 3424
rect 113 3384 115 3464
rect 119 3424 128 3464
rect 119 3384 121 3424
rect 133 3384 135 3424
rect 139 3384 149 3424
rect 153 3384 155 3424
rect 167 3384 169 3424
rect 173 3384 181 3424
rect 185 3384 187 3424
rect 199 3384 201 3424
rect 205 3384 207 3424
rect 245 3384 247 3424
rect 251 3384 255 3424
rect 259 3404 270 3424
rect 296 3404 305 3464
rect 259 3384 261 3404
rect 273 3384 275 3404
rect 279 3384 283 3404
rect 287 3384 291 3404
rect 303 3384 305 3404
rect 309 3384 311 3464
rect 363 3384 365 3424
rect 369 3384 371 3424
rect 423 3384 425 3424
rect 429 3384 431 3424
rect 443 3384 445 3424
rect 449 3384 451 3424
rect 508 3384 510 3424
rect 514 3384 518 3424
rect 530 3384 532 3464
rect 536 3384 540 3464
rect 544 3384 546 3464
rect 608 3384 610 3424
rect 614 3384 618 3424
rect 630 3384 632 3464
rect 636 3384 640 3464
rect 644 3384 646 3464
rect 689 3384 691 3424
rect 695 3384 697 3424
rect 709 3384 711 3424
rect 715 3384 717 3424
rect 769 3384 771 3464
rect 775 3384 781 3464
rect 785 3384 787 3464
rect 809 3384 811 3464
rect 815 3384 821 3464
rect 825 3384 827 3464
rect 1037 3456 1051 3464
rect 889 3384 891 3424
rect 895 3384 897 3424
rect 963 3384 965 3424
rect 969 3420 985 3424
rect 969 3384 971 3420
rect 983 3384 985 3420
rect 989 3384 991 3424
rect 1003 3384 1005 3424
rect 1009 3384 1011 3424
rect 1049 3384 1051 3456
rect 1055 3452 1071 3464
rect 1055 3384 1057 3452
rect 1069 3384 1071 3452
rect 1075 3384 1077 3464
rect 1089 3384 1091 3464
rect 1095 3384 1097 3464
rect 1149 3384 1151 3464
rect 1155 3384 1159 3464
rect 1163 3384 1165 3464
rect 1229 3384 1231 3424
rect 1235 3384 1237 3424
rect 1249 3384 1251 3424
rect 1255 3384 1257 3424
rect 1309 3384 1311 3424
rect 1315 3384 1317 3424
rect 1329 3384 1331 3424
rect 1335 3384 1337 3424
rect 1394 3384 1396 3464
rect 1400 3384 1404 3464
rect 1408 3384 1410 3464
rect 1422 3384 1426 3424
rect 1430 3384 1432 3424
rect 1493 3384 1495 3464
rect 1499 3424 1508 3464
rect 1499 3384 1501 3424
rect 1513 3384 1515 3424
rect 1519 3384 1529 3424
rect 1533 3384 1535 3424
rect 1547 3384 1549 3424
rect 1553 3384 1561 3424
rect 1565 3384 1567 3424
rect 1579 3384 1581 3424
rect 1585 3384 1587 3424
rect 1625 3384 1627 3424
rect 1631 3384 1635 3424
rect 1639 3404 1650 3424
rect 1676 3404 1685 3464
rect 1639 3384 1641 3404
rect 1653 3384 1655 3404
rect 1659 3384 1663 3404
rect 1667 3384 1671 3404
rect 1683 3384 1685 3404
rect 1689 3384 1691 3464
rect 1743 3384 1745 3424
rect 1749 3384 1751 3424
rect 1763 3384 1765 3424
rect 1769 3384 1771 3424
rect 1814 3384 1816 3464
rect 1820 3384 1824 3464
rect 1828 3384 1830 3464
rect 1842 3384 1846 3424
rect 1850 3384 1852 3424
rect 1909 3384 1911 3464
rect 1915 3384 1917 3464
rect 1983 3384 1985 3424
rect 1989 3384 1991 3424
rect 2003 3384 2005 3424
rect 2009 3384 2011 3424
rect 2059 3384 2061 3464
rect 2065 3384 2067 3464
rect 2079 3384 2083 3424
rect 2087 3384 2091 3424
rect 2103 3384 2105 3424
rect 2109 3384 2111 3424
rect 2149 3384 2151 3424
rect 2155 3384 2157 3424
rect 2169 3384 2171 3424
rect 2175 3384 2177 3424
rect 2229 3384 2231 3424
rect 2235 3384 2237 3424
rect 2249 3384 2251 3424
rect 2255 3420 2271 3424
rect 2255 3384 2257 3420
rect 2269 3384 2271 3420
rect 2275 3384 2277 3424
rect 2329 3384 2331 3424
rect 2335 3384 2337 3424
rect 2389 3384 2391 3424
rect 2395 3384 2397 3424
rect 2449 3384 2451 3464
rect 2455 3404 2464 3464
rect 2632 3424 2641 3464
rect 2490 3404 2501 3424
rect 2455 3384 2457 3404
rect 2469 3384 2473 3404
rect 2477 3384 2481 3404
rect 2485 3384 2487 3404
rect 2499 3384 2501 3404
rect 2505 3384 2509 3424
rect 2513 3384 2515 3424
rect 2553 3384 2555 3424
rect 2559 3384 2561 3424
rect 2573 3384 2575 3424
rect 2579 3384 2587 3424
rect 2591 3384 2593 3424
rect 2605 3384 2607 3424
rect 2611 3384 2621 3424
rect 2625 3384 2627 3424
rect 2639 3384 2641 3424
rect 2645 3384 2647 3464
rect 2694 3384 2696 3464
rect 2700 3384 2704 3464
rect 2708 3384 2710 3464
rect 2722 3384 2726 3424
rect 2730 3384 2732 3424
rect 2789 3384 2791 3424
rect 2795 3384 2799 3424
rect 2811 3384 2813 3464
rect 2817 3384 2819 3464
rect 2869 3384 2871 3424
rect 2875 3384 2877 3424
rect 2889 3384 2891 3424
rect 2895 3384 2897 3424
rect 2949 3384 2951 3464
rect 2955 3404 2964 3464
rect 3132 3424 3141 3464
rect 2990 3404 3001 3424
rect 2955 3384 2957 3404
rect 2969 3384 2973 3404
rect 2977 3384 2981 3404
rect 2985 3384 2987 3404
rect 2999 3384 3001 3404
rect 3005 3384 3009 3424
rect 3013 3384 3015 3424
rect 3053 3384 3055 3424
rect 3059 3384 3061 3424
rect 3073 3384 3075 3424
rect 3079 3384 3087 3424
rect 3091 3384 3093 3424
rect 3105 3384 3107 3424
rect 3111 3384 3121 3424
rect 3125 3384 3127 3424
rect 3139 3384 3141 3424
rect 3145 3384 3147 3464
rect 3208 3384 3210 3424
rect 3214 3384 3218 3424
rect 3230 3384 3232 3464
rect 3236 3384 3240 3464
rect 3244 3384 3246 3464
rect 3303 3384 3305 3424
rect 3309 3384 3311 3424
rect 3349 3384 3351 3464
rect 3355 3384 3359 3464
rect 3363 3384 3365 3464
rect 3429 3384 3431 3424
rect 3435 3384 3437 3424
rect 3515 3384 3517 3464
rect 3521 3384 3525 3464
rect 3529 3384 3531 3464
rect 3557 3456 3571 3464
rect 3569 3384 3571 3456
rect 3575 3452 3591 3464
rect 3575 3384 3577 3452
rect 3589 3384 3591 3452
rect 3595 3384 3597 3464
rect 3609 3384 3611 3464
rect 3615 3384 3617 3464
rect 3669 3384 3671 3464
rect 3675 3384 3681 3464
rect 3685 3463 3701 3464
rect 3685 3384 3687 3463
rect 3699 3384 3701 3463
rect 3705 3463 3719 3464
rect 3705 3384 3707 3463
rect 3783 3384 3785 3464
rect 3789 3396 3791 3464
rect 3803 3396 3805 3464
rect 3789 3384 3805 3396
rect 3809 3462 3825 3464
rect 3809 3384 3811 3462
rect 3823 3384 3825 3462
rect 3829 3450 3845 3464
rect 3829 3384 3831 3450
rect 3843 3384 3845 3450
rect 3849 3462 3863 3464
rect 3849 3384 3851 3462
rect 3903 3384 3905 3424
rect 3909 3384 3911 3424
rect 3923 3384 3925 3424
rect 3929 3384 3931 3424
rect 3969 3384 3971 3464
rect 3975 3404 3984 3464
rect 4152 3424 4161 3464
rect 4010 3404 4021 3424
rect 3975 3384 3977 3404
rect 3989 3384 3993 3404
rect 3997 3384 4001 3404
rect 4005 3384 4007 3404
rect 4019 3384 4021 3404
rect 4025 3384 4029 3424
rect 4033 3384 4035 3424
rect 4073 3384 4075 3424
rect 4079 3384 4081 3424
rect 4093 3384 4095 3424
rect 4099 3384 4107 3424
rect 4111 3384 4113 3424
rect 4125 3384 4127 3424
rect 4131 3384 4141 3424
rect 4145 3384 4147 3424
rect 4159 3384 4161 3424
rect 4165 3384 4167 3464
rect 4209 3384 4211 3464
rect 4215 3404 4224 3464
rect 4392 3424 4401 3464
rect 4250 3404 4261 3424
rect 4215 3384 4217 3404
rect 4229 3384 4233 3404
rect 4237 3384 4241 3404
rect 4245 3384 4247 3404
rect 4259 3384 4261 3404
rect 4265 3384 4269 3424
rect 4273 3384 4275 3424
rect 4313 3384 4315 3424
rect 4319 3384 4321 3424
rect 4333 3384 4335 3424
rect 4339 3384 4347 3424
rect 4351 3384 4353 3424
rect 4365 3384 4367 3424
rect 4371 3384 4381 3424
rect 4385 3384 4387 3424
rect 4399 3384 4401 3424
rect 4405 3384 4407 3464
rect 4463 3384 4465 3464
rect 4469 3384 4471 3464
rect 4483 3384 4485 3464
rect 4489 3384 4491 3464
rect 4503 3384 4505 3464
rect 4509 3384 4511 3464
rect 4523 3384 4525 3464
rect 4529 3384 4531 3464
rect 4543 3384 4545 3464
rect 4549 3384 4551 3464
rect 4563 3384 4565 3464
rect 4569 3384 4571 3464
rect 4583 3384 4585 3464
rect 4589 3384 4591 3464
rect 4603 3384 4605 3464
rect 4609 3384 4611 3464
rect 4654 3384 4656 3464
rect 4660 3384 4664 3464
rect 4668 3384 4670 3464
rect 4682 3384 4686 3424
rect 4690 3384 4692 3424
rect 33 3276 35 3356
rect 39 3316 41 3356
rect 53 3316 55 3356
rect 59 3316 69 3356
rect 73 3316 75 3356
rect 87 3316 89 3356
rect 93 3316 101 3356
rect 105 3316 107 3356
rect 119 3316 121 3356
rect 125 3316 127 3356
rect 165 3316 167 3356
rect 171 3316 175 3356
rect 179 3336 181 3356
rect 193 3336 195 3356
rect 199 3336 203 3356
rect 207 3336 211 3356
rect 223 3336 225 3356
rect 179 3316 190 3336
rect 39 3276 48 3316
rect 216 3276 225 3336
rect 229 3276 231 3356
rect 283 3276 285 3356
rect 289 3344 305 3356
rect 289 3276 291 3344
rect 303 3276 305 3344
rect 309 3278 311 3356
rect 323 3278 325 3356
rect 309 3276 325 3278
rect 329 3290 331 3356
rect 343 3290 345 3356
rect 329 3276 345 3290
rect 349 3278 351 3356
rect 403 3316 405 3356
rect 409 3316 411 3356
rect 423 3316 425 3356
rect 429 3316 431 3356
rect 349 3276 363 3278
rect 469 3276 471 3356
rect 475 3336 477 3356
rect 489 3336 493 3356
rect 497 3336 501 3356
rect 505 3336 507 3356
rect 519 3336 521 3356
rect 475 3276 484 3336
rect 510 3316 521 3336
rect 525 3316 529 3356
rect 533 3316 535 3356
rect 573 3316 575 3356
rect 579 3316 581 3356
rect 593 3316 595 3356
rect 599 3316 607 3356
rect 611 3316 613 3356
rect 625 3316 627 3356
rect 631 3316 641 3356
rect 645 3316 647 3356
rect 659 3316 661 3356
rect 652 3276 661 3316
rect 665 3276 667 3356
rect 728 3316 730 3356
rect 734 3316 738 3356
rect 750 3276 752 3356
rect 756 3276 760 3356
rect 764 3276 766 3356
rect 823 3276 825 3356
rect 829 3344 845 3356
rect 829 3276 831 3344
rect 843 3276 845 3344
rect 849 3278 851 3356
rect 863 3278 865 3356
rect 849 3276 865 3278
rect 869 3290 871 3356
rect 883 3290 885 3356
rect 869 3276 885 3290
rect 889 3278 891 3356
rect 929 3316 931 3356
rect 935 3316 937 3356
rect 949 3316 951 3356
rect 955 3316 957 3356
rect 1023 3316 1025 3356
rect 1029 3320 1031 3356
rect 1043 3320 1045 3356
rect 1029 3316 1045 3320
rect 1049 3316 1051 3356
rect 1063 3316 1065 3356
rect 1069 3316 1071 3356
rect 889 3276 903 3278
rect 1119 3276 1121 3356
rect 1125 3276 1127 3356
rect 1139 3316 1143 3356
rect 1147 3316 1151 3356
rect 1163 3316 1165 3356
rect 1169 3316 1171 3356
rect 1209 3316 1211 3356
rect 1215 3316 1217 3356
rect 1229 3316 1231 3356
rect 1235 3320 1237 3356
rect 1249 3320 1251 3356
rect 1235 3316 1251 3320
rect 1255 3316 1257 3356
rect 1314 3276 1316 3356
rect 1320 3276 1324 3356
rect 1328 3276 1330 3356
rect 1342 3316 1346 3356
rect 1350 3316 1352 3356
rect 1409 3316 1411 3356
rect 1415 3316 1417 3356
rect 1429 3316 1431 3356
rect 1435 3316 1437 3356
rect 1513 3277 1515 3356
rect 1501 3276 1515 3277
rect 1519 3277 1521 3356
rect 1533 3277 1535 3356
rect 1519 3276 1535 3277
rect 1539 3276 1545 3356
rect 1549 3276 1551 3356
rect 1603 3316 1605 3356
rect 1609 3316 1611 3356
rect 1623 3316 1625 3356
rect 1629 3316 1631 3356
rect 1674 3276 1676 3356
rect 1680 3276 1684 3356
rect 1688 3276 1690 3356
rect 1702 3316 1706 3356
rect 1710 3316 1712 3356
rect 1788 3316 1790 3356
rect 1794 3316 1798 3356
rect 1810 3276 1812 3356
rect 1816 3276 1820 3356
rect 1824 3276 1826 3356
rect 1869 3316 1871 3356
rect 1875 3316 1877 3356
rect 1889 3316 1891 3356
rect 1895 3316 1897 3356
rect 1954 3276 1956 3356
rect 1960 3276 1964 3356
rect 1968 3276 1970 3356
rect 1982 3316 1986 3356
rect 1990 3316 1992 3356
rect 2068 3316 2070 3356
rect 2074 3316 2078 3356
rect 2090 3276 2092 3356
rect 2096 3276 2100 3356
rect 2104 3276 2106 3356
rect 2149 3316 2151 3356
rect 2155 3316 2157 3356
rect 2214 3276 2216 3356
rect 2220 3276 2224 3356
rect 2228 3276 2230 3356
rect 2242 3316 2246 3356
rect 2250 3316 2252 3356
rect 2323 3316 2325 3356
rect 2329 3316 2331 3356
rect 2369 3316 2371 3356
rect 2375 3316 2377 3356
rect 2389 3316 2391 3356
rect 2395 3316 2397 3356
rect 2449 3276 2451 3356
rect 2455 3336 2457 3356
rect 2469 3336 2473 3356
rect 2477 3336 2481 3356
rect 2485 3336 2487 3356
rect 2499 3336 2501 3356
rect 2455 3276 2464 3336
rect 2490 3316 2501 3336
rect 2505 3316 2509 3356
rect 2513 3316 2515 3356
rect 2553 3316 2555 3356
rect 2559 3316 2561 3356
rect 2573 3316 2575 3356
rect 2579 3316 2587 3356
rect 2591 3316 2593 3356
rect 2605 3316 2607 3356
rect 2611 3316 2621 3356
rect 2625 3316 2627 3356
rect 2639 3316 2641 3356
rect 2632 3276 2641 3316
rect 2645 3276 2647 3356
rect 2689 3316 2691 3356
rect 2695 3316 2699 3356
rect 2711 3276 2713 3356
rect 2717 3276 2719 3356
rect 2769 3276 2771 3356
rect 2775 3336 2777 3356
rect 2789 3336 2793 3356
rect 2797 3336 2801 3356
rect 2805 3336 2807 3356
rect 2819 3336 2821 3356
rect 2775 3276 2784 3336
rect 2810 3316 2821 3336
rect 2825 3316 2829 3356
rect 2833 3316 2835 3356
rect 2873 3316 2875 3356
rect 2879 3316 2881 3356
rect 2893 3316 2895 3356
rect 2899 3316 2907 3356
rect 2911 3316 2913 3356
rect 2925 3316 2927 3356
rect 2931 3316 2941 3356
rect 2945 3316 2947 3356
rect 2959 3316 2961 3356
rect 2952 3276 2961 3316
rect 2965 3276 2967 3356
rect 3028 3316 3030 3356
rect 3034 3316 3038 3356
rect 3050 3276 3052 3356
rect 3056 3276 3060 3356
rect 3064 3276 3066 3356
rect 3128 3316 3130 3356
rect 3134 3316 3138 3356
rect 3150 3276 3152 3356
rect 3156 3276 3160 3356
rect 3164 3276 3166 3356
rect 3214 3276 3216 3356
rect 3220 3276 3224 3356
rect 3228 3276 3230 3356
rect 3242 3316 3246 3356
rect 3250 3316 3252 3356
rect 3328 3316 3330 3356
rect 3334 3316 3338 3356
rect 3350 3276 3352 3356
rect 3356 3276 3360 3356
rect 3364 3276 3366 3356
rect 3414 3276 3416 3356
rect 3420 3276 3424 3356
rect 3428 3276 3430 3356
rect 3442 3316 3446 3356
rect 3450 3316 3452 3356
rect 3509 3316 3511 3356
rect 3515 3316 3517 3356
rect 3529 3316 3531 3356
rect 3535 3316 3537 3356
rect 3589 3316 3591 3356
rect 3595 3316 3597 3356
rect 3609 3316 3611 3356
rect 3615 3316 3617 3356
rect 3669 3316 3671 3356
rect 3675 3316 3677 3356
rect 3689 3316 3691 3356
rect 3695 3316 3697 3356
rect 3749 3316 3751 3356
rect 3755 3316 3757 3356
rect 3769 3316 3771 3356
rect 3775 3316 3777 3356
rect 3829 3316 3831 3356
rect 3835 3316 3839 3356
rect 3851 3276 3853 3356
rect 3857 3276 3859 3356
rect 3923 3316 3925 3356
rect 3929 3316 3931 3356
rect 3943 3316 3945 3356
rect 3949 3316 3951 3356
rect 4015 3276 4017 3356
rect 4021 3276 4025 3356
rect 4029 3276 4031 3356
rect 4069 3316 4071 3356
rect 4075 3316 4079 3356
rect 4091 3276 4093 3356
rect 4097 3276 4099 3356
rect 4163 3316 4165 3356
rect 4169 3316 4171 3356
rect 4228 3316 4230 3356
rect 4234 3316 4238 3356
rect 4250 3276 4252 3356
rect 4256 3276 4260 3356
rect 4264 3276 4266 3356
rect 4323 3316 4325 3356
rect 4329 3316 4331 3356
rect 4374 3276 4376 3356
rect 4380 3276 4384 3356
rect 4388 3276 4390 3356
rect 4402 3316 4406 3356
rect 4410 3316 4412 3356
rect 4483 3316 4485 3356
rect 4489 3316 4491 3356
rect 4503 3316 4505 3356
rect 4509 3316 4511 3356
rect 4553 3276 4555 3356
rect 4559 3316 4561 3356
rect 4573 3316 4575 3356
rect 4579 3316 4589 3356
rect 4593 3316 4595 3356
rect 4607 3316 4609 3356
rect 4613 3316 4621 3356
rect 4625 3316 4627 3356
rect 4639 3316 4641 3356
rect 4645 3316 4647 3356
rect 4685 3316 4687 3356
rect 4691 3316 4695 3356
rect 4699 3336 4701 3356
rect 4713 3336 4715 3356
rect 4719 3336 4723 3356
rect 4727 3336 4731 3356
rect 4743 3336 4745 3356
rect 4699 3316 4710 3336
rect 4559 3276 4568 3316
rect 4736 3276 4745 3336
rect 4749 3276 4751 3356
rect 43 2904 45 2984
rect 49 2916 51 2984
rect 63 2916 65 2984
rect 49 2904 65 2916
rect 69 2982 85 2984
rect 69 2904 71 2982
rect 83 2904 85 2982
rect 89 2970 105 2984
rect 89 2904 91 2970
rect 103 2904 105 2970
rect 109 2982 123 2984
rect 109 2904 111 2982
rect 159 2904 161 2984
rect 165 2904 167 2984
rect 179 2904 183 2944
rect 187 2904 191 2944
rect 203 2904 205 2944
rect 209 2904 211 2944
rect 249 2904 251 2984
rect 255 2924 264 2984
rect 432 2944 441 2984
rect 290 2924 301 2944
rect 255 2904 257 2924
rect 269 2904 273 2924
rect 277 2904 281 2924
rect 285 2904 287 2924
rect 299 2904 301 2924
rect 305 2904 309 2944
rect 313 2904 315 2944
rect 353 2904 355 2944
rect 359 2904 361 2944
rect 373 2904 375 2944
rect 379 2904 387 2944
rect 391 2904 393 2944
rect 405 2904 407 2944
rect 411 2904 421 2944
rect 425 2904 427 2944
rect 439 2904 441 2944
rect 445 2904 447 2984
rect 494 2904 496 2984
rect 500 2904 504 2984
rect 508 2904 510 2984
rect 522 2904 526 2944
rect 530 2904 532 2944
rect 589 2904 591 2944
rect 595 2904 597 2944
rect 609 2904 611 2944
rect 615 2904 617 2944
rect 683 2904 685 2944
rect 689 2904 691 2944
rect 703 2904 705 2944
rect 709 2904 711 2944
rect 775 2904 777 2984
rect 781 2904 785 2984
rect 789 2904 791 2984
rect 829 2904 831 2944
rect 835 2904 837 2944
rect 849 2904 851 2944
rect 855 2904 857 2944
rect 928 2904 930 2944
rect 934 2904 938 2944
rect 950 2904 952 2984
rect 956 2904 960 2984
rect 964 2904 966 2984
rect 1028 2904 1030 2944
rect 1034 2904 1038 2944
rect 1050 2904 1052 2984
rect 1056 2904 1060 2984
rect 1064 2904 1066 2984
rect 1135 2904 1137 2984
rect 1141 2904 1145 2984
rect 1149 2904 1151 2984
rect 1208 2904 1210 2944
rect 1214 2904 1218 2944
rect 1230 2904 1232 2984
rect 1236 2904 1240 2984
rect 1244 2904 1246 2984
rect 1289 2904 1291 2944
rect 1295 2904 1297 2944
rect 1309 2904 1311 2944
rect 1315 2904 1317 2944
rect 1383 2904 1385 2984
rect 1389 2904 1391 2984
rect 1429 2904 1431 2944
rect 1435 2904 1437 2944
rect 1449 2904 1451 2944
rect 1455 2904 1457 2944
rect 1509 2904 1511 2944
rect 1515 2904 1517 2944
rect 1529 2904 1531 2944
rect 1535 2904 1537 2944
rect 1589 2904 1591 2944
rect 1595 2904 1599 2944
rect 1611 2904 1613 2984
rect 1617 2904 1619 2984
rect 1674 2904 1676 2984
rect 1680 2904 1684 2984
rect 1688 2904 1690 2984
rect 1702 2904 1706 2944
rect 1710 2904 1712 2944
rect 1774 2904 1776 2984
rect 1780 2904 1784 2984
rect 1788 2904 1790 2984
rect 1802 2904 1806 2944
rect 1810 2904 1812 2944
rect 1869 2904 1871 2984
rect 1875 2904 1879 2984
rect 1883 2904 1885 2984
rect 1937 2976 1951 2984
rect 1949 2904 1951 2976
rect 1955 2972 1971 2984
rect 1955 2904 1957 2972
rect 1969 2904 1971 2972
rect 1975 2904 1977 2984
rect 1989 2904 1991 2984
rect 1995 2904 1997 2984
rect 2049 2904 2051 2944
rect 2055 2904 2057 2944
rect 2114 2904 2116 2984
rect 2120 2904 2124 2984
rect 2128 2904 2130 2984
rect 2142 2904 2146 2944
rect 2150 2904 2152 2944
rect 2209 2904 2211 2984
rect 2215 2904 2219 2984
rect 2223 2904 2225 2984
rect 2303 2904 2305 2944
rect 2309 2904 2311 2944
rect 2323 2904 2325 2944
rect 2329 2904 2331 2944
rect 2374 2904 2376 2984
rect 2380 2904 2384 2984
rect 2388 2904 2390 2984
rect 2402 2904 2406 2944
rect 2410 2904 2412 2944
rect 2469 2904 2471 2944
rect 2475 2904 2477 2944
rect 2534 2904 2536 2984
rect 2540 2904 2544 2984
rect 2548 2904 2550 2984
rect 2562 2904 2566 2944
rect 2570 2904 2572 2944
rect 2629 2904 2631 2944
rect 2635 2904 2639 2944
rect 2651 2904 2653 2984
rect 2657 2904 2659 2984
rect 2709 2904 2711 2944
rect 2715 2904 2717 2944
rect 2729 2904 2731 2944
rect 2735 2904 2737 2944
rect 2793 2904 2795 2984
rect 2799 2944 2808 2984
rect 2799 2904 2801 2944
rect 2813 2904 2815 2944
rect 2819 2904 2829 2944
rect 2833 2904 2835 2944
rect 2847 2904 2849 2944
rect 2853 2904 2861 2944
rect 2865 2904 2867 2944
rect 2879 2904 2881 2944
rect 2885 2904 2887 2944
rect 2925 2904 2927 2944
rect 2931 2904 2935 2944
rect 2939 2924 2950 2944
rect 2976 2924 2985 2984
rect 2939 2904 2941 2924
rect 2953 2904 2955 2924
rect 2959 2904 2963 2924
rect 2967 2904 2971 2924
rect 2983 2904 2985 2924
rect 2989 2904 2991 2984
rect 3055 2904 3057 2984
rect 3061 2904 3065 2984
rect 3069 2904 3071 2984
rect 3123 2904 3125 2984
rect 3129 2904 3131 2984
rect 3143 2904 3145 2984
rect 3149 2972 3165 2984
rect 3149 2904 3151 2972
rect 3163 2904 3165 2972
rect 3169 2976 3183 2984
rect 3169 2904 3171 2976
rect 3209 2904 3211 2984
rect 3215 2904 3219 2984
rect 3223 2904 3225 2984
rect 3293 2904 3295 2984
rect 3299 2944 3308 2984
rect 3299 2904 3301 2944
rect 3313 2904 3315 2944
rect 3319 2904 3329 2944
rect 3333 2904 3335 2944
rect 3347 2904 3349 2944
rect 3353 2904 3361 2944
rect 3365 2904 3367 2944
rect 3379 2904 3381 2944
rect 3385 2904 3387 2944
rect 3425 2904 3427 2944
rect 3431 2904 3435 2944
rect 3439 2924 3450 2944
rect 3476 2924 3485 2984
rect 3439 2904 3441 2924
rect 3453 2904 3455 2924
rect 3459 2904 3463 2924
rect 3467 2904 3471 2924
rect 3483 2904 3485 2924
rect 3489 2904 3491 2984
rect 3533 2904 3535 2984
rect 3539 2944 3548 2984
rect 3539 2904 3541 2944
rect 3553 2904 3555 2944
rect 3559 2904 3569 2944
rect 3573 2904 3575 2944
rect 3587 2904 3589 2944
rect 3593 2904 3601 2944
rect 3605 2904 3607 2944
rect 3619 2904 3621 2944
rect 3625 2904 3627 2944
rect 3665 2904 3667 2944
rect 3671 2904 3675 2944
rect 3679 2924 3690 2944
rect 3716 2924 3725 2984
rect 3679 2904 3681 2924
rect 3693 2904 3695 2924
rect 3699 2904 3703 2924
rect 3707 2904 3711 2924
rect 3723 2904 3725 2924
rect 3729 2904 3731 2984
rect 3769 2904 3771 2984
rect 3775 2904 3779 2984
rect 3783 2904 3785 2984
rect 3868 2904 3870 2944
rect 3874 2904 3878 2944
rect 3890 2904 3892 2984
rect 3896 2904 3900 2984
rect 3904 2904 3906 2984
rect 3968 2904 3970 2944
rect 3974 2904 3978 2944
rect 3990 2904 3992 2984
rect 3996 2904 4000 2984
rect 4004 2904 4006 2984
rect 4054 2904 4056 2984
rect 4060 2904 4064 2984
rect 4068 2904 4070 2984
rect 4082 2904 4086 2944
rect 4090 2904 4092 2944
rect 4154 2904 4156 2984
rect 4160 2904 4164 2984
rect 4168 2904 4170 2984
rect 4182 2904 4186 2944
rect 4190 2904 4192 2944
rect 4249 2904 4251 2944
rect 4255 2904 4257 2944
rect 4309 2904 4311 2944
rect 4315 2904 4317 2944
rect 4329 2904 4331 2944
rect 4335 2940 4351 2944
rect 4335 2904 4337 2940
rect 4349 2904 4351 2940
rect 4355 2904 4357 2944
rect 4409 2904 4411 2984
rect 4415 2924 4424 2984
rect 4592 2944 4601 2984
rect 4450 2924 4461 2944
rect 4415 2904 4417 2924
rect 4429 2904 4433 2924
rect 4437 2904 4441 2924
rect 4445 2904 4447 2924
rect 4459 2904 4461 2924
rect 4465 2904 4469 2944
rect 4473 2904 4475 2944
rect 4513 2904 4515 2944
rect 4519 2904 4521 2944
rect 4533 2904 4535 2944
rect 4539 2904 4547 2944
rect 4551 2904 4553 2944
rect 4565 2904 4567 2944
rect 4571 2904 4581 2944
rect 4585 2904 4587 2944
rect 4599 2904 4601 2944
rect 4605 2904 4607 2984
rect 4654 2904 4656 2984
rect 4660 2904 4664 2984
rect 4668 2904 4670 2984
rect 4682 2904 4686 2944
rect 4690 2904 4692 2944
rect 43 2836 45 2876
rect 49 2836 51 2876
rect 108 2836 110 2876
rect 114 2836 118 2876
rect 130 2796 132 2876
rect 136 2796 140 2876
rect 144 2796 146 2876
rect 189 2798 191 2876
rect 177 2796 191 2798
rect 195 2810 197 2876
rect 209 2810 211 2876
rect 195 2796 211 2810
rect 215 2798 217 2876
rect 229 2798 231 2876
rect 215 2796 231 2798
rect 235 2864 251 2876
rect 235 2796 237 2864
rect 249 2796 251 2864
rect 255 2796 257 2876
rect 309 2836 311 2876
rect 315 2836 317 2876
rect 329 2836 331 2876
rect 335 2836 337 2876
rect 389 2836 391 2876
rect 395 2836 397 2876
rect 409 2836 413 2876
rect 417 2836 421 2876
rect 433 2796 435 2876
rect 439 2796 441 2876
rect 508 2836 510 2876
rect 514 2836 518 2876
rect 530 2796 532 2876
rect 536 2796 540 2876
rect 544 2796 546 2876
rect 589 2836 591 2876
rect 595 2836 597 2876
rect 609 2836 611 2876
rect 615 2836 617 2876
rect 683 2796 685 2876
rect 689 2796 691 2876
rect 743 2796 745 2876
rect 749 2796 751 2876
rect 789 2836 791 2876
rect 795 2836 797 2876
rect 809 2836 811 2876
rect 815 2836 817 2876
rect 869 2836 871 2876
rect 875 2836 877 2876
rect 889 2836 893 2876
rect 897 2836 901 2876
rect 913 2796 915 2876
rect 919 2796 921 2876
rect 988 2836 990 2876
rect 994 2836 998 2876
rect 1010 2796 1012 2876
rect 1016 2796 1020 2876
rect 1024 2796 1026 2876
rect 1069 2836 1071 2876
rect 1075 2836 1077 2876
rect 1089 2836 1091 2876
rect 1095 2836 1097 2876
rect 1168 2836 1170 2876
rect 1174 2836 1178 2876
rect 1190 2796 1192 2876
rect 1196 2796 1200 2876
rect 1204 2796 1206 2876
rect 1249 2796 1251 2876
rect 1255 2856 1257 2876
rect 1269 2856 1273 2876
rect 1277 2856 1281 2876
rect 1285 2856 1287 2876
rect 1299 2856 1301 2876
rect 1255 2796 1264 2856
rect 1290 2836 1301 2856
rect 1305 2836 1309 2876
rect 1313 2836 1315 2876
rect 1353 2836 1355 2876
rect 1359 2836 1361 2876
rect 1373 2836 1375 2876
rect 1379 2836 1387 2876
rect 1391 2836 1393 2876
rect 1405 2836 1407 2876
rect 1411 2836 1421 2876
rect 1425 2836 1427 2876
rect 1439 2836 1441 2876
rect 1432 2796 1441 2836
rect 1445 2796 1447 2876
rect 1501 2796 1503 2876
rect 1507 2796 1509 2876
rect 1521 2836 1525 2876
rect 1529 2836 1531 2876
rect 1573 2796 1575 2876
rect 1579 2836 1581 2876
rect 1593 2836 1595 2876
rect 1599 2836 1609 2876
rect 1613 2836 1615 2876
rect 1627 2836 1629 2876
rect 1633 2836 1641 2876
rect 1645 2836 1647 2876
rect 1659 2836 1661 2876
rect 1665 2836 1667 2876
rect 1705 2836 1707 2876
rect 1711 2836 1715 2876
rect 1719 2856 1721 2876
rect 1733 2856 1735 2876
rect 1739 2856 1743 2876
rect 1747 2856 1751 2876
rect 1763 2856 1765 2876
rect 1719 2836 1730 2856
rect 1579 2796 1588 2836
rect 1756 2796 1765 2856
rect 1769 2796 1771 2876
rect 1814 2796 1816 2876
rect 1820 2796 1824 2876
rect 1828 2796 1830 2876
rect 1842 2836 1846 2876
rect 1850 2836 1852 2876
rect 1909 2836 1911 2876
rect 1915 2836 1917 2876
rect 1969 2796 1971 2876
rect 1975 2796 1981 2876
rect 1985 2796 1987 2876
rect 2009 2796 2011 2876
rect 2015 2796 2021 2876
rect 2025 2796 2027 2876
rect 2115 2796 2117 2876
rect 2121 2796 2125 2876
rect 2129 2796 2131 2876
rect 2195 2796 2197 2876
rect 2201 2796 2205 2876
rect 2209 2796 2211 2876
rect 2275 2796 2277 2876
rect 2281 2796 2285 2876
rect 2289 2796 2291 2876
rect 2329 2836 2331 2876
rect 2335 2836 2337 2876
rect 2415 2796 2417 2876
rect 2421 2796 2425 2876
rect 2429 2796 2431 2876
rect 2469 2836 2471 2876
rect 2475 2836 2477 2876
rect 2529 2836 2531 2876
rect 2535 2836 2537 2876
rect 2549 2836 2553 2876
rect 2557 2836 2561 2876
rect 2573 2796 2575 2876
rect 2579 2796 2581 2876
rect 2634 2796 2636 2876
rect 2640 2796 2644 2876
rect 2648 2796 2650 2876
rect 2662 2836 2666 2876
rect 2670 2836 2672 2876
rect 2734 2796 2736 2876
rect 2740 2796 2744 2876
rect 2748 2796 2750 2876
rect 2762 2836 2766 2876
rect 2770 2836 2772 2876
rect 2829 2836 2831 2876
rect 2835 2836 2837 2876
rect 2849 2836 2851 2876
rect 2855 2836 2857 2876
rect 2913 2796 2915 2876
rect 2919 2836 2921 2876
rect 2933 2836 2935 2876
rect 2939 2836 2949 2876
rect 2953 2836 2955 2876
rect 2967 2836 2969 2876
rect 2973 2836 2981 2876
rect 2985 2836 2987 2876
rect 2999 2836 3001 2876
rect 3005 2836 3007 2876
rect 3045 2836 3047 2876
rect 3051 2836 3055 2876
rect 3059 2856 3061 2876
rect 3073 2856 3075 2876
rect 3079 2856 3083 2876
rect 3087 2856 3091 2876
rect 3103 2856 3105 2876
rect 3059 2836 3070 2856
rect 2919 2796 2928 2836
rect 3096 2796 3105 2856
rect 3109 2796 3111 2876
rect 3153 2796 3155 2876
rect 3159 2836 3161 2876
rect 3173 2836 3175 2876
rect 3179 2836 3189 2876
rect 3193 2836 3195 2876
rect 3207 2836 3209 2876
rect 3213 2836 3221 2876
rect 3225 2836 3227 2876
rect 3239 2836 3241 2876
rect 3245 2836 3247 2876
rect 3285 2836 3287 2876
rect 3291 2836 3295 2876
rect 3299 2856 3301 2876
rect 3313 2856 3315 2876
rect 3319 2856 3323 2876
rect 3327 2856 3331 2876
rect 3343 2856 3345 2876
rect 3299 2836 3310 2856
rect 3159 2796 3168 2836
rect 3336 2796 3345 2856
rect 3349 2796 3351 2876
rect 3403 2836 3405 2876
rect 3409 2836 3411 2876
rect 3475 2796 3477 2876
rect 3481 2796 3485 2876
rect 3489 2796 3491 2876
rect 3543 2796 3545 2876
rect 3549 2796 3551 2876
rect 3593 2796 3595 2876
rect 3599 2836 3601 2876
rect 3613 2836 3615 2876
rect 3619 2836 3629 2876
rect 3633 2836 3635 2876
rect 3647 2836 3649 2876
rect 3653 2836 3661 2876
rect 3665 2836 3667 2876
rect 3679 2836 3681 2876
rect 3685 2836 3687 2876
rect 3725 2836 3727 2876
rect 3731 2836 3735 2876
rect 3739 2856 3741 2876
rect 3753 2856 3755 2876
rect 3759 2856 3763 2876
rect 3767 2856 3771 2876
rect 3783 2856 3785 2876
rect 3739 2836 3750 2856
rect 3599 2796 3608 2836
rect 3776 2796 3785 2856
rect 3789 2796 3791 2876
rect 3843 2796 3845 2876
rect 3849 2864 3865 2876
rect 3849 2796 3851 2864
rect 3863 2796 3865 2864
rect 3869 2798 3871 2876
rect 3883 2798 3885 2876
rect 3869 2796 3885 2798
rect 3889 2810 3891 2876
rect 3903 2810 3905 2876
rect 3889 2796 3905 2810
rect 3909 2798 3911 2876
rect 3909 2796 3923 2798
rect 3975 2796 3977 2876
rect 3981 2796 3985 2876
rect 3989 2796 3991 2876
rect 4034 2796 4036 2876
rect 4040 2796 4044 2876
rect 4048 2796 4050 2876
rect 4062 2836 4066 2876
rect 4070 2836 4072 2876
rect 4148 2836 4150 2876
rect 4154 2836 4158 2876
rect 4170 2796 4172 2876
rect 4176 2796 4180 2876
rect 4184 2796 4186 2876
rect 4229 2796 4231 2876
rect 4235 2796 4239 2876
rect 4243 2796 4245 2876
rect 4313 2796 4315 2876
rect 4319 2836 4321 2876
rect 4333 2836 4335 2876
rect 4339 2836 4349 2876
rect 4353 2836 4355 2876
rect 4367 2836 4369 2876
rect 4373 2836 4381 2876
rect 4385 2836 4387 2876
rect 4399 2836 4401 2876
rect 4405 2836 4407 2876
rect 4445 2836 4447 2876
rect 4451 2836 4455 2876
rect 4459 2856 4461 2876
rect 4473 2856 4475 2876
rect 4479 2856 4483 2876
rect 4487 2856 4491 2876
rect 4503 2856 4505 2876
rect 4459 2836 4470 2856
rect 4319 2796 4328 2836
rect 4496 2796 4505 2856
rect 4509 2796 4511 2876
rect 4554 2796 4556 2876
rect 4560 2796 4564 2876
rect 4568 2796 4570 2876
rect 4582 2836 4586 2876
rect 4590 2836 4592 2876
rect 4649 2836 4651 2876
rect 4655 2836 4657 2876
rect 4669 2836 4671 2876
rect 4675 2836 4677 2876
rect 117 2496 131 2504
rect 29 2424 31 2464
rect 35 2424 37 2464
rect 49 2424 51 2464
rect 55 2460 71 2464
rect 55 2424 57 2460
rect 69 2424 71 2460
rect 75 2424 77 2464
rect 129 2424 131 2496
rect 135 2492 151 2504
rect 135 2424 137 2492
rect 149 2424 151 2492
rect 155 2424 157 2504
rect 169 2424 171 2504
rect 175 2424 177 2504
rect 243 2424 245 2464
rect 249 2424 251 2464
rect 299 2424 301 2504
rect 305 2424 307 2504
rect 319 2424 323 2464
rect 327 2424 331 2464
rect 343 2424 345 2464
rect 349 2424 351 2464
rect 403 2424 405 2504
rect 409 2424 411 2504
rect 423 2424 425 2504
rect 429 2492 445 2504
rect 429 2424 431 2492
rect 443 2424 445 2492
rect 449 2496 463 2504
rect 449 2424 451 2496
rect 503 2424 505 2464
rect 509 2460 525 2464
rect 509 2424 511 2460
rect 523 2424 525 2460
rect 529 2424 531 2464
rect 543 2424 545 2464
rect 549 2424 551 2464
rect 608 2424 610 2464
rect 614 2424 618 2464
rect 630 2424 632 2504
rect 636 2424 640 2504
rect 644 2424 646 2504
rect 703 2424 705 2504
rect 709 2424 711 2504
rect 763 2424 765 2464
rect 769 2424 771 2464
rect 783 2424 785 2464
rect 789 2424 791 2464
rect 843 2424 845 2464
rect 849 2460 865 2464
rect 849 2424 851 2460
rect 863 2424 865 2460
rect 869 2424 871 2464
rect 883 2424 885 2464
rect 889 2424 891 2464
rect 948 2424 950 2464
rect 954 2424 958 2464
rect 970 2424 972 2504
rect 976 2424 980 2504
rect 984 2424 986 2504
rect 1029 2424 1031 2464
rect 1035 2424 1037 2464
rect 1049 2424 1051 2464
rect 1055 2424 1057 2464
rect 1123 2424 1125 2464
rect 1129 2460 1145 2464
rect 1129 2424 1131 2460
rect 1143 2424 1145 2460
rect 1149 2424 1151 2464
rect 1163 2424 1165 2464
rect 1169 2424 1171 2464
rect 1223 2424 1225 2464
rect 1229 2424 1231 2464
rect 1288 2424 1290 2464
rect 1294 2424 1298 2464
rect 1310 2424 1312 2504
rect 1316 2424 1320 2504
rect 1324 2424 1326 2504
rect 1369 2424 1371 2464
rect 1375 2424 1377 2464
rect 1389 2424 1391 2464
rect 1395 2424 1397 2464
rect 1449 2424 1451 2504
rect 1455 2424 1457 2504
rect 1523 2424 1525 2464
rect 1529 2424 1531 2464
rect 1543 2424 1545 2464
rect 1549 2424 1551 2464
rect 1593 2424 1595 2504
rect 1599 2464 1608 2504
rect 1599 2424 1601 2464
rect 1613 2424 1615 2464
rect 1619 2424 1629 2464
rect 1633 2424 1635 2464
rect 1647 2424 1649 2464
rect 1653 2424 1661 2464
rect 1665 2424 1667 2464
rect 1679 2424 1681 2464
rect 1685 2424 1687 2464
rect 1725 2424 1727 2464
rect 1731 2424 1735 2464
rect 1739 2444 1750 2464
rect 1776 2444 1785 2504
rect 1739 2424 1741 2444
rect 1753 2424 1755 2444
rect 1759 2424 1763 2444
rect 1767 2424 1771 2444
rect 1783 2424 1785 2444
rect 1789 2424 1791 2504
rect 1829 2424 1831 2464
rect 1835 2424 1837 2464
rect 1849 2424 1851 2464
rect 1855 2424 1857 2464
rect 1909 2424 1911 2464
rect 1915 2424 1917 2464
rect 1929 2424 1931 2464
rect 1935 2424 1937 2464
rect 1989 2424 1991 2464
rect 1995 2424 1997 2464
rect 2009 2424 2011 2464
rect 2015 2460 2031 2464
rect 2015 2424 2017 2460
rect 2029 2424 2031 2460
rect 2035 2424 2037 2464
rect 2089 2424 2091 2504
rect 2095 2424 2099 2504
rect 2103 2424 2105 2504
rect 2183 2424 2185 2464
rect 2189 2424 2191 2464
rect 2255 2424 2257 2504
rect 2261 2424 2265 2504
rect 2269 2424 2271 2504
rect 2323 2424 2325 2464
rect 2329 2424 2331 2464
rect 2388 2424 2390 2464
rect 2394 2424 2398 2464
rect 2410 2424 2412 2504
rect 2416 2424 2420 2504
rect 2424 2424 2426 2504
rect 2469 2424 2471 2504
rect 2475 2424 2479 2504
rect 2483 2424 2485 2504
rect 2549 2424 2551 2464
rect 2555 2424 2557 2464
rect 2569 2424 2573 2464
rect 2577 2424 2581 2464
rect 2593 2424 2595 2504
rect 2599 2424 2601 2504
rect 2654 2424 2656 2504
rect 2660 2424 2664 2504
rect 2668 2424 2670 2504
rect 2682 2424 2686 2464
rect 2690 2424 2692 2464
rect 2763 2424 2765 2464
rect 2769 2424 2771 2464
rect 2783 2424 2785 2464
rect 2789 2424 2791 2464
rect 2829 2424 2831 2504
rect 2835 2424 2841 2504
rect 2845 2503 2861 2504
rect 2845 2424 2847 2503
rect 2859 2424 2861 2503
rect 2865 2503 2879 2504
rect 2865 2424 2867 2503
rect 2929 2424 2931 2464
rect 2935 2424 2937 2464
rect 2949 2424 2951 2464
rect 2955 2424 2957 2464
rect 3009 2424 3011 2464
rect 3015 2424 3019 2464
rect 3031 2424 3033 2504
rect 3037 2424 3039 2504
rect 3094 2424 3096 2504
rect 3100 2424 3104 2504
rect 3108 2424 3110 2504
rect 3122 2424 3126 2464
rect 3130 2424 3132 2464
rect 3201 2424 3203 2504
rect 3207 2424 3209 2504
rect 3337 2502 3351 2504
rect 3221 2424 3225 2464
rect 3229 2424 3231 2464
rect 3283 2424 3285 2464
rect 3289 2424 3291 2464
rect 3303 2424 3305 2464
rect 3309 2424 3311 2464
rect 3349 2424 3351 2502
rect 3355 2490 3371 2504
rect 3355 2424 3357 2490
rect 3369 2424 3371 2490
rect 3375 2502 3391 2504
rect 3375 2424 3377 2502
rect 3389 2424 3391 2502
rect 3395 2436 3397 2504
rect 3409 2436 3411 2504
rect 3395 2424 3411 2436
rect 3415 2424 3417 2504
rect 3469 2424 3471 2464
rect 3475 2424 3479 2464
rect 3491 2424 3493 2504
rect 3497 2424 3499 2504
rect 3561 2424 3563 2504
rect 3567 2424 3569 2504
rect 3581 2424 3585 2464
rect 3589 2424 3591 2464
rect 3633 2424 3635 2504
rect 3639 2464 3648 2504
rect 3639 2424 3641 2464
rect 3653 2424 3655 2464
rect 3659 2424 3669 2464
rect 3673 2424 3675 2464
rect 3687 2424 3689 2464
rect 3693 2424 3701 2464
rect 3705 2424 3707 2464
rect 3719 2424 3721 2464
rect 3725 2424 3727 2464
rect 3765 2424 3767 2464
rect 3771 2424 3775 2464
rect 3779 2444 3790 2464
rect 3816 2444 3825 2504
rect 3779 2424 3781 2444
rect 3793 2424 3795 2444
rect 3799 2424 3803 2444
rect 3807 2424 3811 2444
rect 3823 2424 3825 2444
rect 3829 2424 3831 2504
rect 3883 2424 3885 2504
rect 3889 2424 3891 2504
rect 3903 2424 3905 2504
rect 3909 2492 3925 2504
rect 3909 2424 3911 2492
rect 3923 2424 3925 2492
rect 3929 2496 3943 2504
rect 3929 2424 3931 2496
rect 3969 2424 3971 2504
rect 3975 2424 3979 2504
rect 3983 2424 3985 2504
rect 4049 2424 4051 2504
rect 4055 2424 4057 2504
rect 4069 2424 4071 2504
rect 4075 2424 4077 2504
rect 4089 2424 4091 2504
rect 4095 2424 4097 2504
rect 4109 2424 4111 2504
rect 4115 2424 4117 2504
rect 4129 2424 4131 2504
rect 4135 2424 4137 2504
rect 4149 2424 4151 2504
rect 4155 2424 4157 2504
rect 4169 2424 4171 2504
rect 4175 2424 4177 2504
rect 4189 2424 4191 2504
rect 4195 2424 4197 2504
rect 4253 2424 4255 2504
rect 4259 2464 4268 2504
rect 4259 2424 4261 2464
rect 4273 2424 4275 2464
rect 4279 2424 4289 2464
rect 4293 2424 4295 2464
rect 4307 2424 4309 2464
rect 4313 2424 4321 2464
rect 4325 2424 4327 2464
rect 4339 2424 4341 2464
rect 4345 2424 4347 2464
rect 4385 2424 4387 2464
rect 4391 2424 4395 2464
rect 4399 2444 4410 2464
rect 4436 2444 4445 2504
rect 4399 2424 4401 2444
rect 4413 2424 4415 2444
rect 4419 2424 4423 2444
rect 4427 2424 4431 2444
rect 4443 2424 4445 2444
rect 4449 2424 4451 2504
rect 4494 2424 4496 2504
rect 4500 2424 4504 2504
rect 4508 2424 4510 2504
rect 4522 2424 4526 2464
rect 4530 2424 4532 2464
rect 4589 2424 4591 2464
rect 4595 2424 4597 2464
rect 4609 2424 4611 2464
rect 4615 2424 4617 2464
rect 4669 2424 4671 2464
rect 4675 2424 4677 2464
rect 4689 2424 4691 2464
rect 4695 2424 4697 2464
rect 43 2356 45 2396
rect 49 2360 51 2396
rect 63 2360 65 2396
rect 49 2356 65 2360
rect 69 2356 71 2396
rect 83 2356 85 2396
rect 89 2356 91 2396
rect 148 2356 150 2396
rect 154 2356 158 2396
rect 170 2316 172 2396
rect 176 2316 180 2396
rect 184 2316 186 2396
rect 234 2316 236 2396
rect 240 2316 244 2396
rect 248 2316 250 2396
rect 262 2356 266 2396
rect 270 2356 272 2396
rect 329 2356 331 2396
rect 335 2356 337 2396
rect 349 2356 351 2396
rect 355 2360 357 2396
rect 369 2360 371 2396
rect 355 2356 371 2360
rect 375 2356 377 2396
rect 429 2324 431 2396
rect 417 2316 431 2324
rect 435 2328 437 2396
rect 449 2328 451 2396
rect 435 2316 451 2328
rect 455 2316 457 2396
rect 469 2316 471 2396
rect 475 2316 477 2396
rect 534 2316 536 2396
rect 540 2316 544 2396
rect 548 2316 550 2396
rect 562 2356 566 2396
rect 570 2356 572 2396
rect 643 2316 645 2396
rect 649 2316 651 2396
rect 663 2316 665 2396
rect 669 2328 671 2396
rect 683 2328 685 2396
rect 669 2316 685 2328
rect 689 2324 691 2396
rect 729 2356 731 2396
rect 735 2356 737 2396
rect 689 2316 703 2324
rect 799 2316 801 2396
rect 805 2316 807 2396
rect 819 2356 823 2396
rect 827 2356 831 2396
rect 843 2356 845 2396
rect 849 2356 851 2396
rect 889 2356 891 2396
rect 895 2356 897 2396
rect 909 2356 911 2396
rect 915 2356 917 2396
rect 969 2356 971 2396
rect 975 2356 977 2396
rect 989 2356 993 2396
rect 997 2356 1001 2396
rect 1013 2316 1015 2396
rect 1019 2316 1021 2396
rect 1088 2356 1090 2396
rect 1094 2356 1098 2396
rect 1110 2316 1112 2396
rect 1116 2316 1120 2396
rect 1124 2316 1126 2396
rect 1188 2356 1190 2396
rect 1194 2356 1198 2396
rect 1210 2316 1212 2396
rect 1216 2316 1220 2396
rect 1224 2316 1226 2396
rect 1273 2316 1275 2396
rect 1279 2356 1281 2396
rect 1293 2356 1295 2396
rect 1299 2356 1309 2396
rect 1313 2356 1315 2396
rect 1327 2356 1329 2396
rect 1333 2356 1341 2396
rect 1345 2356 1347 2396
rect 1359 2356 1361 2396
rect 1365 2356 1367 2396
rect 1405 2356 1407 2396
rect 1411 2356 1415 2396
rect 1419 2376 1421 2396
rect 1433 2376 1435 2396
rect 1439 2376 1443 2396
rect 1447 2376 1451 2396
rect 1463 2376 1465 2396
rect 1419 2356 1430 2376
rect 1279 2316 1288 2356
rect 1456 2316 1465 2376
rect 1469 2316 1471 2396
rect 1528 2356 1530 2396
rect 1534 2356 1538 2396
rect 1550 2316 1552 2396
rect 1556 2316 1560 2396
rect 1564 2316 1566 2396
rect 1613 2316 1615 2396
rect 1619 2356 1621 2396
rect 1633 2356 1635 2396
rect 1639 2356 1649 2396
rect 1653 2356 1655 2396
rect 1667 2356 1669 2396
rect 1673 2356 1681 2396
rect 1685 2356 1687 2396
rect 1699 2356 1701 2396
rect 1705 2356 1707 2396
rect 1745 2356 1747 2396
rect 1751 2356 1755 2396
rect 1759 2376 1761 2396
rect 1773 2376 1775 2396
rect 1779 2376 1783 2396
rect 1787 2376 1791 2396
rect 1803 2376 1805 2396
rect 1759 2356 1770 2376
rect 1619 2316 1628 2356
rect 1796 2316 1805 2376
rect 1809 2316 1811 2396
rect 1863 2356 1865 2396
rect 1869 2356 1871 2396
rect 1923 2356 1925 2396
rect 1929 2356 1931 2396
rect 1974 2316 1976 2396
rect 1980 2316 1984 2396
rect 1988 2316 1990 2396
rect 2002 2356 2006 2396
rect 2010 2356 2012 2396
rect 2073 2316 2075 2396
rect 2079 2356 2081 2396
rect 2093 2356 2095 2396
rect 2099 2356 2109 2396
rect 2113 2356 2115 2396
rect 2127 2356 2129 2396
rect 2133 2356 2141 2396
rect 2145 2356 2147 2396
rect 2159 2356 2161 2396
rect 2165 2356 2167 2396
rect 2205 2356 2207 2396
rect 2211 2356 2215 2396
rect 2219 2376 2221 2396
rect 2233 2376 2235 2396
rect 2239 2376 2243 2396
rect 2247 2376 2251 2396
rect 2263 2376 2265 2396
rect 2219 2356 2230 2376
rect 2079 2316 2088 2356
rect 2256 2316 2265 2376
rect 2269 2316 2271 2396
rect 2323 2316 2325 2396
rect 2329 2316 2331 2396
rect 2343 2316 2345 2396
rect 2349 2328 2351 2396
rect 2363 2328 2365 2396
rect 2349 2316 2365 2328
rect 2369 2324 2371 2396
rect 2369 2316 2383 2324
rect 2423 2316 2425 2396
rect 2429 2316 2431 2396
rect 2443 2316 2445 2396
rect 2449 2328 2451 2396
rect 2463 2328 2465 2396
rect 2449 2316 2465 2328
rect 2469 2324 2471 2396
rect 2509 2356 2511 2396
rect 2515 2356 2517 2396
rect 2529 2356 2531 2396
rect 2535 2360 2537 2396
rect 2549 2360 2551 2396
rect 2535 2356 2551 2360
rect 2555 2356 2557 2396
rect 2609 2356 2611 2396
rect 2615 2356 2617 2396
rect 2629 2356 2633 2396
rect 2637 2356 2641 2396
rect 2469 2316 2483 2324
rect 2653 2316 2655 2396
rect 2659 2316 2661 2396
rect 2709 2316 2711 2396
rect 2715 2376 2717 2396
rect 2729 2376 2733 2396
rect 2737 2376 2741 2396
rect 2745 2376 2747 2396
rect 2759 2376 2761 2396
rect 2715 2316 2724 2376
rect 2750 2356 2761 2376
rect 2765 2356 2769 2396
rect 2773 2356 2775 2396
rect 2813 2356 2815 2396
rect 2819 2356 2821 2396
rect 2833 2356 2835 2396
rect 2839 2356 2847 2396
rect 2851 2356 2853 2396
rect 2865 2356 2867 2396
rect 2871 2356 2881 2396
rect 2885 2356 2887 2396
rect 2899 2356 2901 2396
rect 2892 2316 2901 2356
rect 2905 2316 2907 2396
rect 2968 2356 2970 2396
rect 2974 2356 2978 2396
rect 2990 2316 2992 2396
rect 2996 2316 3000 2396
rect 3004 2316 3006 2396
rect 3068 2356 3070 2396
rect 3074 2356 3078 2396
rect 3090 2316 3092 2396
rect 3096 2316 3100 2396
rect 3104 2316 3106 2396
rect 3154 2316 3156 2396
rect 3160 2316 3164 2396
rect 3168 2316 3170 2396
rect 3182 2356 3186 2396
rect 3190 2356 3192 2396
rect 3249 2316 3251 2396
rect 3255 2376 3257 2396
rect 3269 2376 3273 2396
rect 3277 2376 3281 2396
rect 3285 2376 3287 2396
rect 3299 2376 3301 2396
rect 3255 2316 3264 2376
rect 3290 2356 3301 2376
rect 3305 2356 3309 2396
rect 3313 2356 3315 2396
rect 3353 2356 3355 2396
rect 3359 2356 3361 2396
rect 3373 2356 3375 2396
rect 3379 2356 3387 2396
rect 3391 2356 3393 2396
rect 3405 2356 3407 2396
rect 3411 2356 3421 2396
rect 3425 2356 3427 2396
rect 3439 2356 3441 2396
rect 3432 2316 3441 2356
rect 3445 2316 3447 2396
rect 3508 2356 3510 2396
rect 3514 2356 3518 2396
rect 3530 2316 3532 2396
rect 3536 2316 3540 2396
rect 3544 2316 3546 2396
rect 3615 2316 3617 2396
rect 3621 2316 3625 2396
rect 3629 2316 3631 2396
rect 3669 2316 3671 2396
rect 3675 2316 3681 2396
rect 3685 2317 3687 2396
rect 3699 2317 3701 2396
rect 3685 2316 3701 2317
rect 3705 2317 3707 2396
rect 3783 2356 3785 2396
rect 3789 2356 3791 2396
rect 3803 2356 3805 2396
rect 3809 2356 3811 2396
rect 3705 2316 3719 2317
rect 3863 2316 3865 2396
rect 3869 2384 3885 2396
rect 3869 2316 3871 2384
rect 3883 2316 3885 2384
rect 3889 2318 3891 2396
rect 3903 2318 3905 2396
rect 3889 2316 3905 2318
rect 3909 2330 3911 2396
rect 3923 2330 3925 2396
rect 3909 2316 3925 2330
rect 3929 2318 3931 2396
rect 3929 2316 3943 2318
rect 3983 2316 3985 2396
rect 3989 2384 4005 2396
rect 3989 2316 3991 2384
rect 4003 2316 4005 2384
rect 4009 2318 4011 2396
rect 4023 2318 4025 2396
rect 4009 2316 4025 2318
rect 4029 2330 4031 2396
rect 4043 2330 4045 2396
rect 4029 2316 4045 2330
rect 4049 2318 4051 2396
rect 4049 2316 4063 2318
rect 4093 2316 4095 2396
rect 4099 2356 4101 2396
rect 4113 2356 4115 2396
rect 4119 2356 4129 2396
rect 4133 2356 4135 2396
rect 4147 2356 4149 2396
rect 4153 2356 4161 2396
rect 4165 2356 4167 2396
rect 4179 2356 4181 2396
rect 4185 2356 4187 2396
rect 4225 2356 4227 2396
rect 4231 2356 4235 2396
rect 4239 2376 4241 2396
rect 4253 2376 4255 2396
rect 4259 2376 4263 2396
rect 4267 2376 4271 2396
rect 4283 2376 4285 2396
rect 4239 2356 4250 2376
rect 4099 2316 4108 2356
rect 4276 2316 4285 2376
rect 4289 2316 4291 2396
rect 4329 2316 4331 2396
rect 4335 2376 4337 2396
rect 4349 2376 4353 2396
rect 4357 2376 4361 2396
rect 4365 2376 4367 2396
rect 4379 2376 4381 2396
rect 4335 2316 4344 2376
rect 4370 2356 4381 2376
rect 4385 2356 4389 2396
rect 4393 2356 4395 2396
rect 4433 2356 4435 2396
rect 4439 2356 4441 2396
rect 4453 2356 4455 2396
rect 4459 2356 4467 2396
rect 4471 2356 4473 2396
rect 4485 2356 4487 2396
rect 4491 2356 4501 2396
rect 4505 2356 4507 2396
rect 4519 2356 4521 2396
rect 4512 2316 4521 2356
rect 4525 2316 4527 2396
rect 4574 2316 4576 2396
rect 4580 2316 4584 2396
rect 4588 2316 4590 2396
rect 4602 2356 4606 2396
rect 4610 2356 4612 2396
rect 4669 2356 4671 2396
rect 4675 2356 4677 2396
rect 4689 2356 4691 2396
rect 4695 2356 4697 2396
rect 41 1944 43 2024
rect 47 1944 49 2024
rect 61 1944 65 1984
rect 69 1944 71 1984
rect 128 1944 130 1984
rect 134 1944 138 1984
rect 150 1944 152 2024
rect 156 1944 160 2024
rect 164 1944 166 2024
rect 297 2016 311 2024
rect 223 1944 225 1984
rect 229 1980 245 1984
rect 229 1944 231 1980
rect 243 1944 245 1980
rect 249 1944 251 1984
rect 263 1944 265 1984
rect 269 1944 271 1984
rect 309 1944 311 2016
rect 315 2012 331 2024
rect 315 1944 317 2012
rect 329 1944 331 2012
rect 335 1944 337 2024
rect 349 1944 351 2024
rect 355 1944 357 2024
rect 397 2016 411 2024
rect 409 1944 411 2016
rect 415 2012 431 2024
rect 415 1944 417 2012
rect 429 1944 431 2012
rect 435 1944 437 2024
rect 449 1944 451 2024
rect 455 1944 457 2024
rect 697 2016 711 2024
rect 509 1944 511 1984
rect 515 1944 517 1984
rect 529 1944 531 1984
rect 535 1980 551 1984
rect 535 1944 537 1980
rect 549 1944 551 1980
rect 555 1944 557 1984
rect 609 1944 611 1984
rect 615 1944 617 1984
rect 629 1944 631 1984
rect 635 1980 651 1984
rect 635 1944 637 1980
rect 649 1944 651 1980
rect 655 1944 657 1984
rect 709 1944 711 2016
rect 715 2012 731 2024
rect 715 1944 717 2012
rect 729 1944 731 2012
rect 735 1944 737 2024
rect 749 1944 751 2024
rect 755 1944 757 2024
rect 828 1944 830 1984
rect 834 1944 838 1984
rect 850 1944 852 2024
rect 856 1944 860 2024
rect 864 1944 866 2024
rect 1197 2016 1211 2024
rect 909 1944 911 1984
rect 915 1944 917 1984
rect 929 1944 931 1984
rect 935 1980 951 1984
rect 935 1944 937 1980
rect 949 1944 951 1980
rect 955 1944 957 1984
rect 1009 1944 1011 1984
rect 1015 1944 1017 1984
rect 1029 1944 1031 1984
rect 1035 1980 1051 1984
rect 1035 1944 1037 1980
rect 1049 1944 1051 1980
rect 1055 1944 1057 1984
rect 1109 1944 1111 1984
rect 1115 1944 1117 1984
rect 1129 1944 1131 1984
rect 1135 1980 1151 1984
rect 1135 1944 1137 1980
rect 1149 1944 1151 1980
rect 1155 1944 1157 1984
rect 1209 1944 1211 2016
rect 1215 2012 1231 2024
rect 1215 1944 1217 2012
rect 1229 1944 1231 2012
rect 1235 1944 1237 2024
rect 1249 1944 1251 2024
rect 1255 1944 1257 2024
rect 1309 1944 1311 2024
rect 1315 1944 1319 2024
rect 1323 1944 1325 2024
rect 1403 1944 1405 1984
rect 1409 1944 1411 1984
rect 1423 1944 1425 1984
rect 1429 1944 1431 1984
rect 1483 1944 1485 1984
rect 1489 1944 1491 1984
rect 1503 1944 1505 1984
rect 1509 1944 1511 1984
rect 1549 1944 1551 1984
rect 1555 1944 1557 1984
rect 1569 1944 1571 1984
rect 1575 1944 1577 1984
rect 1648 1944 1650 1984
rect 1654 1944 1658 1984
rect 1670 1944 1672 2024
rect 1676 1944 1680 2024
rect 1684 1944 1686 2024
rect 1717 2016 1731 2024
rect 1729 1944 1731 2016
rect 1735 2012 1751 2024
rect 1735 1944 1737 2012
rect 1749 1944 1751 2012
rect 1755 1944 1757 2024
rect 1769 1944 1771 2024
rect 1775 1944 1777 2024
rect 1829 1944 1831 2024
rect 1835 1944 1839 2024
rect 1843 1944 1845 2024
rect 1928 1944 1930 1984
rect 1934 1944 1938 1984
rect 1950 1944 1952 2024
rect 1956 1944 1960 2024
rect 1964 1944 1966 2024
rect 2014 1944 2016 2024
rect 2020 1944 2024 2024
rect 2028 1944 2030 2024
rect 2042 1944 2046 1984
rect 2050 1944 2052 1984
rect 2128 1944 2130 1984
rect 2134 1944 2138 1984
rect 2150 1944 2152 2024
rect 2156 1944 2160 2024
rect 2164 1944 2166 2024
rect 2223 1944 2225 2024
rect 2229 1944 2231 2024
rect 2243 1944 2245 2024
rect 2249 1944 2251 2024
rect 2263 1944 2265 2024
rect 2269 1944 2271 2024
rect 2283 1944 2285 2024
rect 2289 1944 2291 2024
rect 2303 1944 2305 2024
rect 2309 1944 2311 2024
rect 2323 1944 2325 2024
rect 2329 1944 2331 2024
rect 2343 1944 2345 2024
rect 2349 1944 2351 2024
rect 2363 1944 2365 2024
rect 2369 1944 2371 2024
rect 2409 1944 2411 1984
rect 2415 1944 2417 1984
rect 2429 1944 2431 1984
rect 2435 1944 2437 1984
rect 2499 1944 2501 2024
rect 2505 1944 2507 2024
rect 2519 1944 2523 1984
rect 2527 1944 2531 1984
rect 2543 1944 2545 1984
rect 2549 1944 2551 1984
rect 2589 1944 2591 2024
rect 2595 1944 2601 2024
rect 2605 2023 2621 2024
rect 2605 1944 2607 2023
rect 2619 1944 2621 2023
rect 2625 2023 2639 2024
rect 2625 1944 2627 2023
rect 2703 1944 2705 1984
rect 2709 1944 2711 1984
rect 2723 1944 2725 1984
rect 2729 1944 2731 1984
rect 2769 1944 2771 1984
rect 2775 1944 2777 1984
rect 2789 1944 2791 1984
rect 2795 1944 2797 1984
rect 2853 1944 2855 2024
rect 2859 1984 2868 2024
rect 2859 1944 2861 1984
rect 2873 1944 2875 1984
rect 2879 1944 2889 1984
rect 2893 1944 2895 1984
rect 2907 1944 2909 1984
rect 2913 1944 2921 1984
rect 2925 1944 2927 1984
rect 2939 1944 2941 1984
rect 2945 1944 2947 1984
rect 2985 1944 2987 1984
rect 2991 1944 2995 1984
rect 2999 1964 3010 1984
rect 3036 1964 3045 2024
rect 2999 1944 3001 1964
rect 3013 1944 3015 1964
rect 3019 1944 3023 1964
rect 3027 1944 3031 1964
rect 3043 1944 3045 1964
rect 3049 1944 3051 2024
rect 3103 1944 3105 2024
rect 3109 1944 3111 2024
rect 3123 1944 3125 2024
rect 3129 2012 3145 2024
rect 3129 1944 3131 2012
rect 3143 1944 3145 2012
rect 3149 2016 3163 2024
rect 3149 1944 3151 2016
rect 3189 1944 3191 2024
rect 3195 1944 3199 2024
rect 3203 1944 3205 2024
rect 3283 1944 3285 2024
rect 3289 1956 3291 2024
rect 3303 1956 3305 2024
rect 3289 1944 3305 1956
rect 3309 2022 3325 2024
rect 3309 1944 3311 2022
rect 3323 1944 3325 2022
rect 3329 2010 3345 2024
rect 3329 1944 3331 2010
rect 3343 1944 3345 2010
rect 3349 2022 3363 2024
rect 3349 1944 3351 2022
rect 3393 1944 3395 2024
rect 3399 1984 3408 2024
rect 3399 1944 3401 1984
rect 3413 1944 3415 1984
rect 3419 1944 3429 1984
rect 3433 1944 3435 1984
rect 3447 1944 3449 1984
rect 3453 1944 3461 1984
rect 3465 1944 3467 1984
rect 3479 1944 3481 1984
rect 3485 1944 3487 1984
rect 3525 1944 3527 1984
rect 3531 1944 3535 1984
rect 3539 1964 3550 1984
rect 3576 1964 3585 2024
rect 3539 1944 3541 1964
rect 3553 1944 3555 1964
rect 3559 1944 3563 1964
rect 3567 1944 3571 1964
rect 3583 1944 3585 1964
rect 3589 1944 3591 2024
rect 3634 1944 3636 2024
rect 3640 1944 3644 2024
rect 3648 1944 3650 2024
rect 3662 1944 3666 1984
rect 3670 1944 3672 1984
rect 3733 1944 3735 2024
rect 3739 1984 3748 2024
rect 3739 1944 3741 1984
rect 3753 1944 3755 1984
rect 3759 1944 3769 1984
rect 3773 1944 3775 1984
rect 3787 1944 3789 1984
rect 3793 1944 3801 1984
rect 3805 1944 3807 1984
rect 3819 1944 3821 1984
rect 3825 1944 3827 1984
rect 3865 1944 3867 1984
rect 3871 1944 3875 1984
rect 3879 1964 3890 1984
rect 3916 1964 3925 2024
rect 3879 1944 3881 1964
rect 3893 1944 3895 1964
rect 3899 1944 3903 1964
rect 3907 1944 3911 1964
rect 3923 1944 3925 1964
rect 3929 1944 3931 2024
rect 3969 1944 3971 2024
rect 3975 1964 3984 2024
rect 4152 1984 4161 2024
rect 4010 1964 4021 1984
rect 3975 1944 3977 1964
rect 3989 1944 3993 1964
rect 3997 1944 4001 1964
rect 4005 1944 4007 1964
rect 4019 1944 4021 1964
rect 4025 1944 4029 1984
rect 4033 1944 4035 1984
rect 4073 1944 4075 1984
rect 4079 1944 4081 1984
rect 4093 1944 4095 1984
rect 4099 1944 4107 1984
rect 4111 1944 4113 1984
rect 4125 1944 4127 1984
rect 4131 1944 4141 1984
rect 4145 1944 4147 1984
rect 4159 1944 4161 1984
rect 4165 1944 4167 2024
rect 4223 1944 4225 2024
rect 4229 1956 4231 2024
rect 4243 1956 4245 2024
rect 4229 1944 4245 1956
rect 4249 2022 4265 2024
rect 4249 1944 4251 2022
rect 4263 1944 4265 2022
rect 4269 2010 4285 2024
rect 4269 1944 4271 2010
rect 4283 1944 4285 2010
rect 4289 2022 4303 2024
rect 4289 1944 4291 2022
rect 4329 1944 4331 1984
rect 4335 1944 4337 1984
rect 4415 1944 4417 2024
rect 4421 1944 4425 2024
rect 4429 1944 4431 2024
rect 4495 1944 4497 2024
rect 4501 1944 4505 2024
rect 4509 1944 4511 2024
rect 4549 1944 4551 2024
rect 4555 1964 4564 2024
rect 4732 1984 4741 2024
rect 4590 1964 4601 1984
rect 4555 1944 4557 1964
rect 4569 1944 4573 1964
rect 4577 1944 4581 1964
rect 4585 1944 4587 1964
rect 4599 1944 4601 1964
rect 4605 1944 4609 1984
rect 4613 1944 4615 1984
rect 4653 1944 4655 1984
rect 4659 1944 4661 1984
rect 4673 1944 4675 1984
rect 4679 1944 4687 1984
rect 4691 1944 4693 1984
rect 4705 1944 4707 1984
rect 4711 1944 4721 1984
rect 4725 1944 4727 1984
rect 4739 1944 4741 1984
rect 4745 1944 4747 2024
rect 43 1836 45 1916
rect 49 1904 65 1916
rect 49 1836 51 1904
rect 63 1836 65 1904
rect 69 1838 71 1916
rect 83 1838 85 1916
rect 69 1836 85 1838
rect 89 1850 91 1916
rect 103 1850 105 1916
rect 89 1836 105 1850
rect 109 1838 111 1916
rect 109 1836 123 1838
rect 154 1836 156 1916
rect 160 1836 164 1916
rect 168 1836 170 1916
rect 182 1876 186 1916
rect 190 1876 192 1916
rect 249 1876 251 1916
rect 255 1876 257 1916
rect 269 1876 271 1916
rect 275 1876 277 1916
rect 343 1876 345 1916
rect 349 1880 351 1916
rect 363 1880 365 1916
rect 349 1876 365 1880
rect 369 1876 371 1916
rect 383 1876 385 1916
rect 389 1876 391 1916
rect 429 1838 431 1916
rect 417 1836 431 1838
rect 435 1850 437 1916
rect 449 1850 451 1916
rect 435 1836 451 1850
rect 455 1838 457 1916
rect 469 1838 471 1916
rect 455 1836 471 1838
rect 475 1904 491 1916
rect 475 1836 477 1904
rect 489 1836 491 1904
rect 495 1836 497 1916
rect 549 1876 551 1916
rect 555 1876 557 1916
rect 569 1876 573 1916
rect 577 1876 581 1916
rect 593 1836 595 1916
rect 599 1836 601 1916
rect 663 1836 665 1916
rect 669 1836 671 1916
rect 709 1876 711 1916
rect 715 1876 719 1916
rect 731 1836 733 1916
rect 737 1836 739 1916
rect 808 1876 810 1916
rect 814 1876 818 1916
rect 830 1836 832 1916
rect 836 1836 840 1916
rect 844 1836 846 1916
rect 894 1836 896 1916
rect 900 1836 904 1916
rect 908 1836 910 1916
rect 922 1876 926 1916
rect 930 1876 932 1916
rect 989 1876 991 1916
rect 995 1876 997 1916
rect 1009 1876 1011 1916
rect 1015 1880 1017 1916
rect 1029 1880 1031 1916
rect 1015 1876 1031 1880
rect 1035 1876 1037 1916
rect 1089 1876 1091 1916
rect 1095 1876 1097 1916
rect 1149 1876 1151 1916
rect 1155 1876 1157 1916
rect 1169 1876 1171 1916
rect 1175 1880 1177 1916
rect 1189 1880 1191 1916
rect 1175 1876 1191 1880
rect 1195 1876 1197 1916
rect 1249 1876 1251 1916
rect 1255 1876 1257 1916
rect 1269 1876 1271 1916
rect 1275 1880 1277 1916
rect 1289 1880 1291 1916
rect 1275 1876 1291 1880
rect 1295 1876 1297 1916
rect 1363 1876 1365 1916
rect 1369 1876 1371 1916
rect 1423 1836 1425 1916
rect 1429 1904 1445 1916
rect 1429 1836 1431 1904
rect 1443 1836 1445 1904
rect 1449 1838 1451 1916
rect 1463 1838 1465 1916
rect 1449 1836 1465 1838
rect 1469 1850 1471 1916
rect 1483 1850 1485 1916
rect 1469 1836 1485 1850
rect 1489 1838 1491 1916
rect 1529 1876 1531 1916
rect 1535 1876 1537 1916
rect 1549 1876 1551 1916
rect 1555 1880 1557 1916
rect 1569 1880 1571 1916
rect 1555 1876 1571 1880
rect 1575 1876 1577 1916
rect 1629 1876 1631 1916
rect 1635 1876 1637 1916
rect 1489 1836 1503 1838
rect 1703 1836 1705 1916
rect 1709 1836 1711 1916
rect 1763 1876 1765 1916
rect 1769 1880 1771 1916
rect 1783 1880 1785 1916
rect 1769 1876 1785 1880
rect 1789 1876 1791 1916
rect 1803 1876 1805 1916
rect 1809 1876 1811 1916
rect 1849 1876 1851 1916
rect 1855 1876 1857 1916
rect 1869 1876 1873 1916
rect 1877 1876 1881 1916
rect 1893 1836 1895 1916
rect 1899 1836 1901 1916
rect 1953 1836 1955 1916
rect 1959 1876 1961 1916
rect 1973 1876 1975 1916
rect 1979 1876 1989 1916
rect 1993 1876 1995 1916
rect 2007 1876 2009 1916
rect 2013 1876 2021 1916
rect 2025 1876 2027 1916
rect 2039 1876 2041 1916
rect 2045 1876 2047 1916
rect 2085 1876 2087 1916
rect 2091 1876 2095 1916
rect 2099 1896 2101 1916
rect 2113 1896 2115 1916
rect 2119 1896 2123 1916
rect 2127 1896 2131 1916
rect 2143 1896 2145 1916
rect 2099 1876 2110 1896
rect 1959 1836 1968 1876
rect 2136 1836 2145 1896
rect 2149 1836 2151 1916
rect 2215 1836 2217 1916
rect 2221 1836 2225 1916
rect 2229 1836 2231 1916
rect 2269 1876 2271 1916
rect 2275 1876 2277 1916
rect 2334 1836 2336 1916
rect 2340 1836 2344 1916
rect 2348 1836 2350 1916
rect 2362 1876 2366 1916
rect 2370 1876 2372 1916
rect 2429 1836 2431 1916
rect 2435 1836 2439 1916
rect 2443 1836 2445 1916
rect 2509 1836 2511 1916
rect 2515 1836 2519 1916
rect 2523 1836 2525 1916
rect 2594 1836 2596 1916
rect 2600 1836 2604 1916
rect 2608 1836 2610 1916
rect 2622 1876 2626 1916
rect 2630 1876 2632 1916
rect 2703 1876 2705 1916
rect 2709 1876 2711 1916
rect 2723 1876 2725 1916
rect 2729 1876 2731 1916
rect 2795 1836 2797 1916
rect 2801 1836 2805 1916
rect 2809 1836 2811 1916
rect 2854 1836 2856 1916
rect 2860 1836 2864 1916
rect 2868 1836 2870 1916
rect 2882 1876 2886 1916
rect 2890 1876 2892 1916
rect 2949 1876 2951 1916
rect 2955 1876 2957 1916
rect 3035 1836 3037 1916
rect 3041 1836 3045 1916
rect 3049 1836 3051 1916
rect 3089 1836 3091 1916
rect 3095 1896 3097 1916
rect 3109 1896 3113 1916
rect 3117 1896 3121 1916
rect 3125 1896 3127 1916
rect 3139 1896 3141 1916
rect 3095 1836 3104 1896
rect 3130 1876 3141 1896
rect 3145 1876 3149 1916
rect 3153 1876 3155 1916
rect 3193 1876 3195 1916
rect 3199 1876 3201 1916
rect 3213 1876 3215 1916
rect 3219 1876 3227 1916
rect 3231 1876 3233 1916
rect 3245 1876 3247 1916
rect 3251 1876 3261 1916
rect 3265 1876 3267 1916
rect 3279 1876 3281 1916
rect 3272 1836 3281 1876
rect 3285 1836 3287 1916
rect 3334 1836 3336 1916
rect 3340 1836 3344 1916
rect 3348 1836 3350 1916
rect 3362 1876 3366 1916
rect 3370 1876 3372 1916
rect 3429 1876 3431 1916
rect 3435 1876 3437 1916
rect 3449 1876 3451 1916
rect 3455 1876 3457 1916
rect 3509 1836 3511 1916
rect 3515 1896 3517 1916
rect 3529 1896 3533 1916
rect 3537 1896 3541 1916
rect 3545 1896 3547 1916
rect 3559 1896 3561 1916
rect 3515 1836 3524 1896
rect 3550 1876 3561 1896
rect 3565 1876 3569 1916
rect 3573 1876 3575 1916
rect 3613 1876 3615 1916
rect 3619 1876 3621 1916
rect 3633 1876 3635 1916
rect 3639 1876 3647 1916
rect 3651 1876 3653 1916
rect 3665 1876 3667 1916
rect 3671 1876 3681 1916
rect 3685 1876 3687 1916
rect 3699 1876 3701 1916
rect 3692 1836 3701 1876
rect 3705 1836 3707 1916
rect 3749 1876 3751 1916
rect 3755 1876 3759 1916
rect 3771 1836 3773 1916
rect 3777 1836 3779 1916
rect 3843 1876 3845 1916
rect 3849 1876 3851 1916
rect 3863 1876 3865 1916
rect 3869 1876 3871 1916
rect 3928 1876 3930 1916
rect 3934 1876 3938 1916
rect 3950 1836 3952 1916
rect 3956 1836 3960 1916
rect 3964 1836 3966 1916
rect 4028 1876 4030 1916
rect 4034 1876 4038 1916
rect 4050 1836 4052 1916
rect 4056 1836 4060 1916
rect 4064 1836 4066 1916
rect 4109 1836 4111 1916
rect 4115 1836 4121 1916
rect 4125 1837 4127 1916
rect 4139 1837 4141 1916
rect 4125 1836 4141 1837
rect 4145 1837 4147 1916
rect 4223 1876 4225 1916
rect 4229 1876 4231 1916
rect 4145 1836 4159 1837
rect 4269 1844 4271 1916
rect 4257 1836 4271 1844
rect 4275 1848 4277 1916
rect 4289 1848 4291 1916
rect 4275 1836 4291 1848
rect 4295 1836 4297 1916
rect 4309 1836 4311 1916
rect 4315 1836 4317 1916
rect 4395 1836 4397 1916
rect 4401 1836 4405 1916
rect 4409 1836 4411 1916
rect 4449 1836 4451 1916
rect 4455 1896 4457 1916
rect 4469 1896 4473 1916
rect 4477 1896 4481 1916
rect 4485 1896 4487 1916
rect 4499 1896 4501 1916
rect 4455 1836 4464 1896
rect 4490 1876 4501 1896
rect 4505 1876 4509 1916
rect 4513 1876 4515 1916
rect 4553 1876 4555 1916
rect 4559 1876 4561 1916
rect 4573 1876 4575 1916
rect 4579 1876 4587 1916
rect 4591 1876 4593 1916
rect 4605 1876 4607 1916
rect 4611 1876 4621 1916
rect 4625 1876 4627 1916
rect 4639 1876 4641 1916
rect 4632 1836 4641 1876
rect 4645 1836 4647 1916
rect 4703 1876 4705 1916
rect 4709 1876 4711 1916
rect 4723 1876 4725 1916
rect 4729 1876 4731 1916
rect 43 1464 45 1504
rect 49 1464 51 1504
rect 103 1464 105 1544
rect 109 1464 111 1544
rect 123 1464 125 1544
rect 129 1532 145 1544
rect 129 1464 131 1532
rect 143 1464 145 1532
rect 149 1536 163 1544
rect 149 1464 151 1536
rect 189 1464 191 1504
rect 195 1464 197 1504
rect 209 1464 211 1504
rect 215 1500 231 1504
rect 215 1464 217 1500
rect 229 1464 231 1500
rect 235 1464 237 1504
rect 289 1464 291 1504
rect 295 1464 297 1504
rect 309 1464 311 1504
rect 315 1464 317 1504
rect 388 1464 390 1504
rect 394 1464 398 1504
rect 410 1464 412 1544
rect 416 1464 420 1544
rect 424 1464 426 1544
rect 481 1464 483 1544
rect 487 1464 489 1544
rect 697 1536 711 1544
rect 501 1464 505 1504
rect 509 1464 511 1504
rect 563 1464 565 1504
rect 569 1464 571 1504
rect 609 1464 611 1504
rect 615 1464 617 1504
rect 629 1464 631 1504
rect 635 1500 651 1504
rect 635 1464 637 1500
rect 649 1464 651 1500
rect 655 1464 657 1504
rect 709 1464 711 1536
rect 715 1532 731 1544
rect 715 1464 717 1532
rect 729 1464 731 1532
rect 735 1464 737 1544
rect 749 1464 751 1544
rect 755 1464 757 1544
rect 897 1536 911 1544
rect 809 1464 811 1504
rect 815 1464 817 1504
rect 829 1464 831 1504
rect 835 1500 851 1504
rect 835 1464 837 1500
rect 849 1464 851 1500
rect 855 1464 857 1504
rect 909 1464 911 1536
rect 915 1532 931 1544
rect 915 1464 917 1532
rect 929 1464 931 1532
rect 935 1464 937 1544
rect 949 1464 951 1544
rect 955 1464 957 1544
rect 1009 1464 1011 1504
rect 1015 1464 1017 1504
rect 1029 1464 1031 1504
rect 1035 1500 1051 1504
rect 1035 1464 1037 1500
rect 1049 1464 1051 1500
rect 1055 1464 1057 1504
rect 1128 1464 1130 1504
rect 1134 1464 1138 1504
rect 1150 1464 1152 1544
rect 1156 1464 1160 1544
rect 1164 1464 1166 1544
rect 1297 1536 1311 1544
rect 1209 1464 1211 1504
rect 1215 1464 1217 1504
rect 1229 1464 1231 1504
rect 1235 1500 1251 1504
rect 1235 1464 1237 1500
rect 1249 1464 1251 1500
rect 1255 1464 1257 1504
rect 1309 1464 1311 1536
rect 1315 1532 1331 1544
rect 1315 1464 1317 1532
rect 1329 1464 1331 1532
rect 1335 1464 1337 1544
rect 1349 1464 1351 1544
rect 1355 1464 1357 1544
rect 1557 1536 1571 1544
rect 1423 1464 1425 1504
rect 1429 1464 1431 1504
rect 1469 1464 1471 1504
rect 1475 1464 1477 1504
rect 1489 1464 1491 1504
rect 1495 1500 1511 1504
rect 1495 1464 1497 1500
rect 1509 1464 1511 1500
rect 1515 1464 1517 1504
rect 1569 1464 1571 1536
rect 1575 1532 1591 1544
rect 1575 1464 1577 1532
rect 1589 1464 1591 1532
rect 1595 1464 1597 1544
rect 1609 1464 1611 1544
rect 1615 1464 1617 1544
rect 1669 1464 1671 1504
rect 1675 1464 1677 1504
rect 1689 1464 1691 1504
rect 1695 1500 1711 1504
rect 1695 1464 1697 1500
rect 1709 1464 1711 1500
rect 1715 1464 1717 1504
rect 1774 1464 1776 1544
rect 1780 1464 1784 1544
rect 1788 1464 1790 1544
rect 1802 1464 1806 1504
rect 1810 1464 1812 1504
rect 1883 1464 1885 1544
rect 1889 1464 1891 1544
rect 1903 1464 1905 1544
rect 1909 1532 1925 1544
rect 1909 1464 1911 1532
rect 1923 1464 1925 1532
rect 1929 1536 1943 1544
rect 1929 1464 1931 1536
rect 1969 1464 1971 1504
rect 1975 1464 1977 1504
rect 2029 1464 2031 1504
rect 2035 1464 2037 1504
rect 2049 1464 2051 1504
rect 2055 1500 2071 1504
rect 2055 1464 2057 1500
rect 2069 1464 2071 1500
rect 2075 1464 2077 1504
rect 2148 1464 2150 1504
rect 2154 1464 2158 1504
rect 2170 1464 2172 1544
rect 2176 1464 2180 1544
rect 2184 1464 2186 1544
rect 2229 1464 2231 1504
rect 2235 1464 2237 1504
rect 2289 1464 2291 1544
rect 2295 1484 2304 1544
rect 2472 1504 2481 1544
rect 2330 1484 2341 1504
rect 2295 1464 2297 1484
rect 2309 1464 2313 1484
rect 2317 1464 2321 1484
rect 2325 1464 2327 1484
rect 2339 1464 2341 1484
rect 2345 1464 2349 1504
rect 2353 1464 2355 1504
rect 2393 1464 2395 1504
rect 2399 1464 2401 1504
rect 2413 1464 2415 1504
rect 2419 1464 2427 1504
rect 2431 1464 2433 1504
rect 2445 1464 2447 1504
rect 2451 1464 2461 1504
rect 2465 1464 2467 1504
rect 2479 1464 2481 1504
rect 2485 1464 2487 1544
rect 2548 1464 2550 1504
rect 2554 1464 2558 1504
rect 2570 1464 2572 1544
rect 2576 1464 2580 1544
rect 2584 1464 2586 1544
rect 2639 1464 2641 1544
rect 2645 1464 2647 1544
rect 2659 1464 2663 1504
rect 2667 1464 2671 1504
rect 2683 1464 2685 1504
rect 2689 1464 2691 1504
rect 2729 1464 2731 1544
rect 2735 1464 2739 1544
rect 2743 1464 2745 1544
rect 2797 1536 2811 1544
rect 2809 1464 2811 1536
rect 2815 1532 2831 1544
rect 2815 1464 2817 1532
rect 2829 1464 2831 1532
rect 2835 1464 2837 1544
rect 2849 1464 2851 1544
rect 2855 1464 2857 1544
rect 2935 1464 2937 1544
rect 2941 1464 2945 1544
rect 2949 1464 2951 1544
rect 3003 1464 3005 1504
rect 3009 1464 3011 1504
rect 3063 1464 3065 1504
rect 3069 1464 3071 1504
rect 3114 1464 3116 1544
rect 3120 1464 3124 1544
rect 3128 1464 3130 1544
rect 3142 1464 3146 1504
rect 3150 1464 3152 1504
rect 3209 1464 3211 1504
rect 3215 1464 3217 1504
rect 3229 1464 3231 1504
rect 3235 1464 3237 1504
rect 3303 1464 3305 1504
rect 3309 1464 3311 1504
rect 3323 1464 3325 1504
rect 3329 1464 3331 1504
rect 3388 1464 3390 1504
rect 3394 1464 3398 1504
rect 3410 1464 3412 1544
rect 3416 1464 3420 1544
rect 3424 1464 3426 1544
rect 3473 1464 3475 1544
rect 3479 1504 3488 1544
rect 3479 1464 3481 1504
rect 3493 1464 3495 1504
rect 3499 1464 3509 1504
rect 3513 1464 3515 1504
rect 3527 1464 3529 1504
rect 3533 1464 3541 1504
rect 3545 1464 3547 1504
rect 3559 1464 3561 1504
rect 3565 1464 3567 1504
rect 3605 1464 3607 1504
rect 3611 1464 3615 1504
rect 3619 1484 3630 1504
rect 3656 1484 3665 1544
rect 3619 1464 3621 1484
rect 3633 1464 3635 1484
rect 3639 1464 3643 1484
rect 3647 1464 3651 1484
rect 3663 1464 3665 1484
rect 3669 1464 3671 1544
rect 3709 1464 3711 1504
rect 3715 1464 3717 1504
rect 3783 1464 3785 1504
rect 3789 1464 3791 1504
rect 3848 1464 3850 1504
rect 3854 1464 3858 1504
rect 3870 1464 3872 1544
rect 3876 1464 3880 1544
rect 3884 1464 3886 1544
rect 3929 1464 3931 1544
rect 3935 1464 3939 1544
rect 3943 1464 3945 1544
rect 4009 1464 4011 1544
rect 4015 1464 4019 1544
rect 4023 1464 4025 1544
rect 4137 1536 4151 1544
rect 4089 1464 4091 1504
rect 4095 1464 4097 1504
rect 4149 1464 4151 1536
rect 4155 1532 4171 1544
rect 4155 1464 4157 1532
rect 4169 1464 4171 1532
rect 4175 1464 4177 1544
rect 4189 1464 4191 1544
rect 4195 1464 4197 1544
rect 4249 1464 4251 1544
rect 4255 1464 4259 1544
rect 4263 1464 4265 1544
rect 4317 1536 4331 1544
rect 4329 1464 4331 1536
rect 4335 1532 4351 1544
rect 4335 1464 4337 1532
rect 4349 1464 4351 1532
rect 4355 1464 4357 1544
rect 4369 1464 4371 1544
rect 4375 1464 4377 1544
rect 4429 1464 4431 1504
rect 4435 1464 4437 1504
rect 4489 1464 4491 1504
rect 4495 1464 4497 1504
rect 4563 1464 4565 1504
rect 4569 1464 4571 1504
rect 4614 1464 4616 1544
rect 4620 1464 4624 1544
rect 4628 1464 4630 1544
rect 4642 1464 4646 1504
rect 4650 1464 4652 1504
rect 4709 1464 4711 1504
rect 4715 1464 4717 1504
rect 4729 1464 4731 1504
rect 4735 1464 4737 1504
rect 43 1356 45 1436
rect 49 1356 51 1436
rect 63 1356 65 1436
rect 69 1368 71 1436
rect 83 1368 85 1436
rect 69 1356 85 1368
rect 89 1364 91 1436
rect 129 1396 131 1436
rect 135 1396 137 1436
rect 149 1396 151 1436
rect 155 1400 157 1436
rect 169 1400 171 1436
rect 155 1396 171 1400
rect 175 1396 177 1436
rect 229 1396 231 1436
rect 235 1396 237 1436
rect 249 1396 251 1436
rect 255 1400 257 1436
rect 269 1400 271 1436
rect 255 1396 271 1400
rect 275 1396 277 1436
rect 343 1396 345 1436
rect 349 1396 351 1436
rect 363 1396 365 1436
rect 369 1396 371 1436
rect 89 1356 103 1364
rect 414 1356 416 1436
rect 420 1356 424 1436
rect 428 1356 430 1436
rect 442 1396 446 1436
rect 450 1396 452 1436
rect 509 1364 511 1436
rect 497 1356 511 1364
rect 515 1368 517 1436
rect 529 1368 531 1436
rect 515 1356 531 1368
rect 535 1356 537 1436
rect 549 1356 551 1436
rect 555 1356 557 1436
rect 614 1356 616 1436
rect 620 1356 624 1436
rect 628 1356 630 1436
rect 642 1396 646 1436
rect 650 1396 652 1436
rect 714 1356 716 1436
rect 720 1356 724 1436
rect 728 1356 730 1436
rect 742 1396 746 1436
rect 750 1396 752 1436
rect 809 1396 811 1436
rect 815 1396 817 1436
rect 829 1396 833 1436
rect 837 1396 841 1436
rect 853 1356 855 1436
rect 859 1356 861 1436
rect 923 1396 925 1436
rect 929 1396 931 1436
rect 943 1396 945 1436
rect 949 1396 951 1436
rect 989 1396 991 1436
rect 995 1396 997 1436
rect 1009 1396 1011 1436
rect 1015 1396 1017 1436
rect 1083 1396 1085 1436
rect 1089 1400 1091 1436
rect 1103 1400 1105 1436
rect 1089 1396 1105 1400
rect 1109 1396 1111 1436
rect 1123 1396 1125 1436
rect 1129 1396 1131 1436
rect 1183 1396 1185 1436
rect 1189 1396 1191 1436
rect 1239 1356 1241 1436
rect 1245 1356 1247 1436
rect 1259 1396 1263 1436
rect 1267 1396 1271 1436
rect 1283 1396 1285 1436
rect 1289 1396 1291 1436
rect 1334 1356 1336 1436
rect 1340 1356 1344 1436
rect 1348 1356 1350 1436
rect 1362 1396 1366 1436
rect 1370 1396 1372 1436
rect 1448 1396 1450 1436
rect 1454 1396 1458 1436
rect 1470 1356 1472 1436
rect 1476 1356 1480 1436
rect 1484 1356 1486 1436
rect 1529 1396 1531 1436
rect 1535 1396 1537 1436
rect 1549 1396 1551 1436
rect 1555 1396 1557 1436
rect 1614 1356 1616 1436
rect 1620 1356 1624 1436
rect 1628 1356 1630 1436
rect 1642 1396 1646 1436
rect 1650 1396 1652 1436
rect 1709 1396 1711 1436
rect 1715 1396 1717 1436
rect 1729 1396 1731 1436
rect 1735 1396 1737 1436
rect 1789 1364 1791 1436
rect 1777 1356 1791 1364
rect 1795 1368 1797 1436
rect 1809 1368 1811 1436
rect 1795 1356 1811 1368
rect 1815 1356 1817 1436
rect 1829 1356 1831 1436
rect 1835 1356 1837 1436
rect 1889 1396 1891 1436
rect 1895 1396 1897 1436
rect 1909 1396 1911 1436
rect 1915 1400 1917 1436
rect 1929 1400 1931 1436
rect 1915 1396 1931 1400
rect 1935 1396 1937 1436
rect 1994 1356 1996 1436
rect 2000 1356 2004 1436
rect 2008 1356 2010 1436
rect 2022 1396 2026 1436
rect 2030 1396 2032 1436
rect 2089 1396 2091 1436
rect 2095 1396 2097 1436
rect 2149 1396 2151 1436
rect 2155 1396 2157 1436
rect 2169 1396 2171 1436
rect 2175 1400 2177 1436
rect 2189 1400 2191 1436
rect 2175 1396 2191 1400
rect 2195 1396 2197 1436
rect 2249 1396 2251 1436
rect 2255 1396 2257 1436
rect 2269 1396 2271 1436
rect 2275 1396 2277 1436
rect 2329 1356 2331 1436
rect 2335 1356 2341 1436
rect 2345 1357 2347 1436
rect 2359 1357 2361 1436
rect 2345 1356 2361 1357
rect 2365 1357 2367 1436
rect 2443 1396 2445 1436
rect 2449 1396 2451 1436
rect 2463 1396 2465 1436
rect 2469 1396 2471 1436
rect 2509 1396 2511 1436
rect 2515 1396 2517 1436
rect 2365 1356 2379 1357
rect 2581 1356 2583 1436
rect 2587 1356 2589 1436
rect 2601 1396 2605 1436
rect 2609 1396 2611 1436
rect 2654 1356 2656 1436
rect 2660 1356 2664 1436
rect 2668 1356 2670 1436
rect 2682 1396 2686 1436
rect 2690 1396 2692 1436
rect 2773 1356 2775 1436
rect 2779 1356 2785 1436
rect 2789 1356 2791 1436
rect 2813 1356 2815 1436
rect 2819 1356 2825 1436
rect 2829 1356 2831 1436
rect 2873 1356 2875 1436
rect 2879 1396 2881 1436
rect 2893 1396 2895 1436
rect 2899 1396 2909 1436
rect 2913 1396 2915 1436
rect 2927 1396 2929 1436
rect 2933 1396 2941 1436
rect 2945 1396 2947 1436
rect 2959 1396 2961 1436
rect 2965 1396 2967 1436
rect 3005 1396 3007 1436
rect 3011 1396 3015 1436
rect 3019 1416 3021 1436
rect 3033 1416 3035 1436
rect 3039 1416 3043 1436
rect 3047 1416 3051 1436
rect 3063 1416 3065 1436
rect 3019 1396 3030 1416
rect 2879 1356 2888 1396
rect 3056 1356 3065 1416
rect 3069 1356 3071 1436
rect 3135 1356 3137 1436
rect 3141 1356 3145 1436
rect 3149 1356 3151 1436
rect 3203 1356 3205 1436
rect 3209 1356 3211 1436
rect 3223 1356 3225 1436
rect 3229 1368 3231 1436
rect 3243 1368 3245 1436
rect 3229 1356 3245 1368
rect 3249 1364 3251 1436
rect 3249 1356 3263 1364
rect 3293 1356 3295 1436
rect 3299 1396 3301 1436
rect 3313 1396 3315 1436
rect 3319 1396 3329 1436
rect 3333 1396 3335 1436
rect 3347 1396 3349 1436
rect 3353 1396 3361 1436
rect 3365 1396 3367 1436
rect 3379 1396 3381 1436
rect 3385 1396 3387 1436
rect 3425 1396 3427 1436
rect 3431 1396 3435 1436
rect 3439 1416 3441 1436
rect 3453 1416 3455 1436
rect 3459 1416 3463 1436
rect 3467 1416 3471 1436
rect 3483 1416 3485 1436
rect 3439 1396 3450 1416
rect 3299 1356 3308 1396
rect 3476 1356 3485 1416
rect 3489 1356 3491 1436
rect 3543 1396 3545 1436
rect 3549 1396 3551 1436
rect 3615 1356 3617 1436
rect 3621 1356 3625 1436
rect 3629 1356 3631 1436
rect 3695 1356 3697 1436
rect 3701 1356 3705 1436
rect 3709 1356 3711 1436
rect 3749 1396 3751 1436
rect 3755 1396 3757 1436
rect 3809 1356 3811 1436
rect 3815 1416 3817 1436
rect 3829 1416 3833 1436
rect 3837 1416 3841 1436
rect 3845 1416 3847 1436
rect 3859 1416 3861 1436
rect 3815 1356 3824 1416
rect 3850 1396 3861 1416
rect 3865 1396 3869 1436
rect 3873 1396 3875 1436
rect 3913 1396 3915 1436
rect 3919 1396 3921 1436
rect 3933 1396 3935 1436
rect 3939 1396 3947 1436
rect 3951 1396 3953 1436
rect 3965 1396 3967 1436
rect 3971 1396 3981 1436
rect 3985 1396 3987 1436
rect 3999 1396 4001 1436
rect 3992 1356 4001 1396
rect 4005 1356 4007 1436
rect 4054 1356 4056 1436
rect 4060 1356 4064 1436
rect 4068 1356 4070 1436
rect 4082 1396 4086 1436
rect 4090 1396 4092 1436
rect 4149 1396 4151 1436
rect 4155 1396 4157 1436
rect 4169 1396 4171 1436
rect 4175 1396 4177 1436
rect 4241 1356 4243 1436
rect 4247 1356 4249 1436
rect 4261 1396 4265 1436
rect 4269 1396 4271 1436
rect 4323 1396 4325 1436
rect 4329 1396 4331 1436
rect 4343 1396 4345 1436
rect 4349 1396 4351 1436
rect 4408 1396 4410 1436
rect 4414 1396 4418 1436
rect 4430 1356 4432 1436
rect 4436 1356 4440 1436
rect 4444 1356 4446 1436
rect 4508 1396 4510 1436
rect 4514 1396 4518 1436
rect 4530 1356 4532 1436
rect 4536 1356 4540 1436
rect 4544 1356 4546 1436
rect 4589 1356 4591 1436
rect 4595 1356 4599 1436
rect 4603 1356 4605 1436
rect 4669 1396 4671 1436
rect 4675 1396 4677 1436
rect 4743 1396 4745 1436
rect 4749 1396 4751 1436
rect 48 984 50 1024
rect 54 984 58 1024
rect 70 984 72 1064
rect 76 984 80 1064
rect 84 984 86 1064
rect 134 984 136 1064
rect 140 984 144 1064
rect 148 984 150 1064
rect 317 1056 331 1064
rect 162 984 166 1024
rect 170 984 172 1024
rect 229 984 231 1024
rect 235 984 237 1024
rect 249 984 251 1024
rect 255 1020 271 1024
rect 255 984 257 1020
rect 269 984 271 1020
rect 275 984 277 1024
rect 329 984 331 1056
rect 335 1052 351 1064
rect 335 984 337 1052
rect 349 984 351 1052
rect 355 984 357 1064
rect 369 984 371 1064
rect 375 984 377 1064
rect 517 1056 531 1064
rect 429 984 431 1024
rect 435 984 437 1024
rect 449 984 451 1024
rect 455 1020 471 1024
rect 455 984 457 1020
rect 469 984 471 1020
rect 475 984 477 1024
rect 529 984 531 1056
rect 535 1052 551 1064
rect 535 984 537 1052
rect 549 984 551 1052
rect 555 984 557 1064
rect 569 984 571 1064
rect 575 984 577 1064
rect 643 984 645 1024
rect 649 984 651 1024
rect 663 984 665 1024
rect 669 984 671 1024
rect 719 984 721 1064
rect 725 984 727 1064
rect 739 984 743 1024
rect 747 984 751 1024
rect 763 984 765 1024
rect 769 984 771 1024
rect 823 984 825 1024
rect 829 1020 845 1024
rect 829 984 831 1020
rect 843 984 845 1020
rect 849 984 851 1024
rect 863 984 865 1024
rect 869 984 871 1024
rect 928 984 930 1024
rect 934 984 938 1024
rect 950 984 952 1064
rect 956 984 960 1064
rect 964 984 966 1064
rect 1014 984 1016 1064
rect 1020 984 1024 1064
rect 1028 984 1030 1064
rect 1042 984 1046 1024
rect 1050 984 1052 1024
rect 1128 984 1130 1024
rect 1134 984 1138 1024
rect 1150 984 1152 1064
rect 1156 984 1160 1064
rect 1164 984 1166 1064
rect 1223 984 1225 1024
rect 1229 984 1231 1024
rect 1243 984 1245 1024
rect 1249 984 1251 1024
rect 1299 984 1301 1064
rect 1305 984 1307 1064
rect 1319 984 1323 1024
rect 1327 984 1331 1024
rect 1343 984 1345 1024
rect 1349 984 1351 1024
rect 1389 984 1391 1024
rect 1395 984 1397 1024
rect 1409 984 1411 1024
rect 1415 984 1417 1024
rect 1483 984 1485 1064
rect 1489 984 1491 1064
rect 1543 984 1545 1024
rect 1549 984 1551 1024
rect 1563 984 1565 1024
rect 1569 984 1571 1024
rect 1623 984 1625 1024
rect 1629 984 1631 1024
rect 1643 984 1645 1024
rect 1649 984 1651 1024
rect 1689 984 1691 1024
rect 1695 984 1697 1024
rect 1709 984 1711 1024
rect 1715 1020 1731 1024
rect 1715 984 1717 1020
rect 1729 984 1731 1020
rect 1735 984 1737 1024
rect 1803 984 1805 1024
rect 1809 984 1811 1024
rect 1823 984 1825 1024
rect 1829 984 1831 1024
rect 1869 984 1871 1024
rect 1875 984 1877 1024
rect 1889 984 1891 1024
rect 1895 1020 1911 1024
rect 1895 984 1897 1020
rect 1909 984 1911 1020
rect 1915 984 1917 1024
rect 1969 984 1971 1024
rect 1975 984 1977 1024
rect 1989 984 1991 1024
rect 1995 984 1997 1024
rect 2063 984 2065 1064
rect 2069 996 2071 1064
rect 2083 996 2085 1064
rect 2069 984 2085 996
rect 2089 1062 2105 1064
rect 2089 984 2091 1062
rect 2103 984 2105 1062
rect 2109 1050 2125 1064
rect 2109 984 2111 1050
rect 2123 984 2125 1050
rect 2129 1062 2143 1064
rect 2129 984 2131 1062
rect 2337 1056 2351 1064
rect 2183 984 2185 1024
rect 2189 1020 2205 1024
rect 2189 984 2191 1020
rect 2203 984 2205 1020
rect 2209 984 2211 1024
rect 2223 984 2225 1024
rect 2229 984 2231 1024
rect 2283 984 2285 1024
rect 2289 984 2291 1024
rect 2303 984 2305 1024
rect 2309 984 2311 1024
rect 2349 984 2351 1056
rect 2355 1052 2371 1064
rect 2355 984 2357 1052
rect 2369 984 2371 1052
rect 2375 984 2377 1064
rect 2389 984 2391 1064
rect 2395 984 2397 1064
rect 2463 984 2465 1024
rect 2469 984 2471 1024
rect 2523 984 2525 1024
rect 2529 984 2531 1024
rect 2543 984 2545 1024
rect 2549 984 2551 1024
rect 2613 984 2615 1064
rect 2619 984 2625 1064
rect 2629 984 2631 1064
rect 2653 984 2655 1064
rect 2659 984 2665 1064
rect 2669 984 2671 1064
rect 2709 984 2711 1024
rect 2715 984 2719 1024
rect 2731 984 2733 1064
rect 2737 984 2739 1064
rect 2793 984 2795 1064
rect 2799 1024 2808 1064
rect 2799 984 2801 1024
rect 2813 984 2815 1024
rect 2819 984 2829 1024
rect 2833 984 2835 1024
rect 2847 984 2849 1024
rect 2853 984 2861 1024
rect 2865 984 2867 1024
rect 2879 984 2881 1024
rect 2885 984 2887 1024
rect 2925 984 2927 1024
rect 2931 984 2935 1024
rect 2939 1004 2950 1024
rect 2976 1004 2985 1064
rect 2939 984 2941 1004
rect 2953 984 2955 1004
rect 2959 984 2963 1004
rect 2967 984 2971 1004
rect 2983 984 2985 1004
rect 2989 984 2991 1064
rect 3029 984 3031 1024
rect 3035 984 3037 1024
rect 3049 984 3051 1024
rect 3055 984 3057 1024
rect 3128 984 3130 1024
rect 3134 984 3138 1024
rect 3150 984 3152 1064
rect 3156 984 3160 1064
rect 3164 984 3166 1064
rect 3209 984 3211 1064
rect 3215 984 3217 1064
rect 3229 984 3231 1064
rect 3235 984 3237 1064
rect 3249 984 3251 1064
rect 3255 984 3257 1064
rect 3269 984 3271 1064
rect 3275 984 3277 1064
rect 3341 984 3343 1064
rect 3347 984 3349 1064
rect 3361 984 3365 1024
rect 3369 984 3371 1024
rect 3409 984 3411 1024
rect 3415 984 3419 1024
rect 3431 984 3433 1064
rect 3437 984 3439 1064
rect 3489 984 3491 1064
rect 3495 984 3497 1064
rect 3509 984 3511 1064
rect 3515 984 3517 1064
rect 3529 984 3531 1064
rect 3535 984 3537 1064
rect 3549 984 3551 1064
rect 3555 984 3557 1064
rect 3569 984 3571 1064
rect 3575 984 3577 1064
rect 3589 984 3591 1064
rect 3595 984 3597 1064
rect 3609 984 3611 1064
rect 3615 984 3617 1064
rect 3629 984 3631 1064
rect 3635 984 3637 1064
rect 3689 984 3691 1064
rect 3695 984 3697 1064
rect 3709 984 3711 1064
rect 3715 984 3717 1064
rect 3729 984 3731 1064
rect 3735 984 3737 1064
rect 3749 984 3751 1064
rect 3755 984 3757 1064
rect 3769 984 3771 1064
rect 3775 984 3777 1064
rect 3789 984 3791 1064
rect 3795 984 3797 1064
rect 3809 984 3811 1064
rect 3815 984 3817 1064
rect 3829 984 3831 1064
rect 3835 984 3837 1064
rect 3889 984 3891 1024
rect 3895 984 3899 1024
rect 3911 984 3913 1064
rect 3917 984 3919 1064
rect 3969 984 3971 1024
rect 3975 984 3977 1024
rect 3989 984 3991 1024
rect 3995 984 3997 1024
rect 4049 984 4051 1064
rect 4055 1004 4064 1064
rect 4232 1024 4241 1064
rect 4090 1004 4101 1024
rect 4055 984 4057 1004
rect 4069 984 4073 1004
rect 4077 984 4081 1004
rect 4085 984 4087 1004
rect 4099 984 4101 1004
rect 4105 984 4109 1024
rect 4113 984 4115 1024
rect 4153 984 4155 1024
rect 4159 984 4161 1024
rect 4173 984 4175 1024
rect 4179 984 4187 1024
rect 4191 984 4193 1024
rect 4205 984 4207 1024
rect 4211 984 4221 1024
rect 4225 984 4227 1024
rect 4239 984 4241 1024
rect 4245 984 4247 1064
rect 4289 984 4291 1024
rect 4295 984 4297 1024
rect 4309 984 4311 1024
rect 4315 984 4317 1024
rect 4374 984 4376 1064
rect 4380 984 4384 1064
rect 4388 984 4390 1064
rect 4402 984 4406 1024
rect 4410 984 4412 1024
rect 4483 984 4485 1024
rect 4489 984 4491 1024
rect 4503 984 4505 1024
rect 4509 984 4511 1024
rect 4554 984 4556 1064
rect 4560 984 4564 1064
rect 4568 984 4570 1064
rect 4582 984 4586 1024
rect 4590 984 4592 1024
rect 4649 984 4651 1024
rect 4655 984 4657 1024
rect 4669 984 4671 1024
rect 4675 1020 4691 1024
rect 4675 984 4677 1020
rect 4689 984 4691 1020
rect 4695 984 4697 1024
rect 43 916 45 956
rect 49 916 51 956
rect 63 916 65 956
rect 69 916 71 956
rect 119 876 121 956
rect 125 876 127 956
rect 139 916 143 956
rect 147 916 151 956
rect 163 916 165 956
rect 169 916 171 956
rect 228 916 230 956
rect 234 916 238 956
rect 250 876 252 956
rect 256 876 260 956
rect 264 876 266 956
rect 323 876 325 956
rect 329 944 345 956
rect 329 876 331 944
rect 343 876 345 944
rect 349 878 351 956
rect 363 878 365 956
rect 349 876 365 878
rect 369 890 371 956
rect 383 890 385 956
rect 369 876 385 890
rect 389 878 391 956
rect 389 876 403 878
rect 441 876 443 956
rect 447 876 449 956
rect 461 916 465 956
rect 469 916 471 956
rect 509 916 511 956
rect 515 916 517 956
rect 583 916 585 956
rect 589 916 591 956
rect 643 876 645 956
rect 649 876 651 956
rect 663 876 665 956
rect 669 888 671 956
rect 683 888 685 956
rect 669 876 685 888
rect 689 884 691 956
rect 729 916 731 956
rect 735 916 737 956
rect 749 916 751 956
rect 755 920 757 956
rect 769 920 771 956
rect 755 916 771 920
rect 775 916 777 956
rect 689 876 703 884
rect 839 876 841 956
rect 845 876 847 956
rect 859 916 863 956
rect 867 916 871 956
rect 883 916 885 956
rect 889 916 891 956
rect 929 916 931 956
rect 935 916 937 956
rect 949 916 951 956
rect 955 916 957 956
rect 1023 916 1025 956
rect 1029 920 1031 956
rect 1043 920 1045 956
rect 1029 916 1045 920
rect 1049 916 1051 956
rect 1063 916 1065 956
rect 1069 916 1071 956
rect 1114 876 1116 956
rect 1120 876 1124 956
rect 1128 876 1130 956
rect 1142 916 1146 956
rect 1150 916 1152 956
rect 1223 916 1225 956
rect 1229 920 1231 956
rect 1243 920 1245 956
rect 1229 916 1245 920
rect 1249 916 1251 956
rect 1263 916 1265 956
rect 1269 916 1271 956
rect 1309 916 1311 956
rect 1315 916 1317 956
rect 1374 876 1376 956
rect 1380 876 1384 956
rect 1388 876 1390 956
rect 1402 916 1406 956
rect 1410 916 1412 956
rect 1483 916 1485 956
rect 1489 916 1491 956
rect 1503 916 1505 956
rect 1509 916 1511 956
rect 1549 916 1551 956
rect 1555 916 1557 956
rect 1569 916 1571 956
rect 1575 916 1577 956
rect 1648 916 1650 956
rect 1654 916 1658 956
rect 1670 876 1672 956
rect 1676 876 1680 956
rect 1684 876 1686 956
rect 1729 916 1731 956
rect 1735 916 1737 956
rect 1749 916 1753 956
rect 1757 916 1761 956
rect 1773 876 1775 956
rect 1779 876 1781 956
rect 1843 916 1845 956
rect 1849 916 1851 956
rect 1903 916 1905 956
rect 1909 916 1911 956
rect 1923 916 1925 956
rect 1929 916 1931 956
rect 1969 916 1971 956
rect 1975 916 1977 956
rect 2043 916 2045 956
rect 2049 920 2051 956
rect 2063 920 2065 956
rect 2049 916 2065 920
rect 2069 916 2071 956
rect 2083 916 2085 956
rect 2089 916 2091 956
rect 2129 916 2131 956
rect 2135 916 2137 956
rect 2194 876 2196 956
rect 2200 876 2204 956
rect 2208 876 2210 956
rect 2222 916 2226 956
rect 2230 916 2232 956
rect 2303 876 2305 956
rect 2309 876 2311 956
rect 2323 876 2325 956
rect 2329 888 2331 956
rect 2343 888 2345 956
rect 2329 876 2345 888
rect 2349 884 2351 956
rect 2389 916 2391 956
rect 2395 916 2397 956
rect 2449 916 2451 956
rect 2455 916 2457 956
rect 2469 916 2471 956
rect 2475 920 2477 956
rect 2489 920 2491 956
rect 2475 916 2491 920
rect 2495 916 2497 956
rect 2563 916 2565 956
rect 2569 920 2571 956
rect 2583 920 2585 956
rect 2569 916 2585 920
rect 2589 916 2591 956
rect 2603 916 2605 956
rect 2609 916 2611 956
rect 2349 876 2363 884
rect 2649 884 2651 956
rect 2637 876 2651 884
rect 2655 888 2657 956
rect 2669 888 2671 956
rect 2655 876 2671 888
rect 2675 876 2677 956
rect 2689 876 2691 956
rect 2695 876 2697 956
rect 2763 916 2765 956
rect 2769 916 2771 956
rect 2783 916 2785 956
rect 2789 916 2791 956
rect 2853 876 2855 956
rect 2859 876 2865 956
rect 2869 876 2871 956
rect 2893 876 2895 956
rect 2899 876 2905 956
rect 2909 876 2911 956
rect 2963 916 2965 956
rect 2969 916 2971 956
rect 3035 876 3037 956
rect 3041 876 3045 956
rect 3049 876 3051 956
rect 3115 876 3117 956
rect 3121 876 3125 956
rect 3129 876 3131 956
rect 3169 916 3171 956
rect 3175 916 3177 956
rect 3234 876 3236 956
rect 3240 876 3244 956
rect 3248 876 3250 956
rect 3262 916 3266 956
rect 3270 916 3272 956
rect 3329 916 3331 956
rect 3335 916 3337 956
rect 3349 916 3351 956
rect 3355 916 3357 956
rect 3409 876 3411 956
rect 3415 936 3417 956
rect 3429 936 3433 956
rect 3437 936 3441 956
rect 3445 936 3447 956
rect 3459 936 3461 956
rect 3415 876 3424 936
rect 3450 916 3461 936
rect 3465 916 3469 956
rect 3473 916 3475 956
rect 3513 916 3515 956
rect 3519 916 3521 956
rect 3533 916 3535 956
rect 3539 916 3547 956
rect 3551 916 3553 956
rect 3565 916 3567 956
rect 3571 916 3581 956
rect 3585 916 3587 956
rect 3599 916 3601 956
rect 3592 876 3601 916
rect 3605 876 3607 956
rect 3649 916 3651 956
rect 3655 916 3659 956
rect 3671 876 3673 956
rect 3677 876 3679 956
rect 3733 876 3735 956
rect 3739 916 3741 956
rect 3753 916 3755 956
rect 3759 916 3769 956
rect 3773 916 3775 956
rect 3787 916 3789 956
rect 3793 916 3801 956
rect 3805 916 3807 956
rect 3819 916 3821 956
rect 3825 916 3827 956
rect 3865 916 3867 956
rect 3871 916 3875 956
rect 3879 936 3881 956
rect 3893 936 3895 956
rect 3899 936 3903 956
rect 3907 936 3911 956
rect 3923 936 3925 956
rect 3879 916 3890 936
rect 3739 876 3748 916
rect 3916 876 3925 936
rect 3929 876 3931 956
rect 3988 916 3990 956
rect 3994 916 3998 956
rect 4010 876 4012 956
rect 4016 876 4020 956
rect 4024 876 4026 956
rect 4069 876 4071 956
rect 4075 936 4077 956
rect 4089 936 4093 956
rect 4097 936 4101 956
rect 4105 936 4107 956
rect 4119 936 4121 956
rect 4075 876 4084 936
rect 4110 916 4121 936
rect 4125 916 4129 956
rect 4133 916 4135 956
rect 4173 916 4175 956
rect 4179 916 4181 956
rect 4193 916 4195 956
rect 4199 916 4207 956
rect 4211 916 4213 956
rect 4225 916 4227 956
rect 4231 916 4241 956
rect 4245 916 4247 956
rect 4259 916 4261 956
rect 4252 876 4261 916
rect 4265 876 4267 956
rect 4313 876 4315 956
rect 4319 916 4321 956
rect 4333 916 4335 956
rect 4339 916 4349 956
rect 4353 916 4355 956
rect 4367 916 4369 956
rect 4373 916 4381 956
rect 4385 916 4387 956
rect 4399 916 4401 956
rect 4405 916 4407 956
rect 4445 916 4447 956
rect 4451 916 4455 956
rect 4459 936 4461 956
rect 4473 936 4475 956
rect 4479 936 4483 956
rect 4487 936 4491 956
rect 4503 936 4505 956
rect 4459 916 4470 936
rect 4319 876 4328 916
rect 4496 876 4505 936
rect 4509 876 4511 956
rect 4554 876 4556 956
rect 4560 876 4564 956
rect 4568 876 4570 956
rect 4582 916 4586 956
rect 4590 916 4592 956
rect 4654 876 4656 956
rect 4660 876 4664 956
rect 4668 876 4670 956
rect 4682 916 4686 956
rect 4690 916 4692 956
rect 55 504 57 584
rect 61 504 65 584
rect 69 504 71 584
rect 123 504 125 584
rect 129 504 131 584
rect 143 504 145 584
rect 149 572 165 584
rect 149 504 151 572
rect 163 504 165 572
rect 169 576 183 584
rect 169 504 171 576
rect 209 504 211 544
rect 215 504 217 544
rect 283 504 285 584
rect 289 504 291 584
rect 303 504 305 584
rect 309 572 325 584
rect 309 504 311 572
rect 323 504 325 572
rect 329 576 343 584
rect 329 504 331 576
rect 369 504 371 544
rect 375 504 377 544
rect 389 504 391 544
rect 395 540 411 544
rect 395 504 397 540
rect 409 504 411 540
rect 415 504 417 544
rect 488 504 490 544
rect 494 504 498 544
rect 510 504 512 584
rect 516 504 520 584
rect 524 504 526 584
rect 581 504 583 584
rect 587 504 589 584
rect 601 504 605 544
rect 609 504 611 544
rect 668 504 670 544
rect 674 504 678 544
rect 690 504 692 584
rect 696 504 700 584
rect 704 504 706 584
rect 761 504 763 584
rect 767 504 769 584
rect 781 504 785 544
rect 789 504 791 544
rect 829 504 831 544
rect 835 504 837 544
rect 849 504 853 544
rect 857 504 861 544
rect 873 504 875 584
rect 879 504 881 584
rect 934 504 936 584
rect 940 504 944 584
rect 948 504 950 584
rect 962 504 966 544
rect 970 504 972 544
rect 1048 504 1050 544
rect 1054 504 1058 544
rect 1070 504 1072 584
rect 1076 504 1080 584
rect 1084 504 1086 584
rect 1143 504 1145 584
rect 1149 504 1151 584
rect 1177 576 1191 584
rect 1189 504 1191 576
rect 1195 572 1211 584
rect 1195 504 1197 572
rect 1209 504 1211 572
rect 1215 504 1217 584
rect 1229 504 1231 584
rect 1235 504 1237 584
rect 1303 504 1305 544
rect 1309 504 1311 544
rect 1354 504 1356 584
rect 1360 504 1364 584
rect 1368 504 1370 584
rect 1382 504 1386 544
rect 1390 504 1392 544
rect 1454 504 1456 584
rect 1460 504 1464 584
rect 1468 504 1470 584
rect 1482 504 1486 544
rect 1490 504 1492 544
rect 1563 504 1565 584
rect 1569 504 1571 584
rect 1583 504 1585 584
rect 1589 572 1605 584
rect 1589 504 1591 572
rect 1603 504 1605 572
rect 1609 576 1623 584
rect 1609 504 1611 576
rect 1637 576 1651 584
rect 1649 504 1651 576
rect 1655 572 1671 584
rect 1655 504 1657 572
rect 1669 504 1671 572
rect 1675 504 1677 584
rect 1689 504 1691 584
rect 1695 504 1697 584
rect 1749 504 1751 544
rect 1755 504 1757 544
rect 1769 504 1771 544
rect 1775 540 1791 544
rect 1775 504 1777 540
rect 1789 504 1791 540
rect 1795 504 1797 544
rect 1854 504 1856 584
rect 1860 504 1864 584
rect 1868 504 1870 584
rect 1882 504 1886 544
rect 1890 504 1892 544
rect 1963 504 1965 584
rect 1969 504 1971 584
rect 1983 504 1985 584
rect 1989 572 2005 584
rect 1989 504 1991 572
rect 2003 504 2005 572
rect 2009 576 2023 584
rect 2009 504 2011 576
rect 2054 504 2056 584
rect 2060 504 2064 584
rect 2068 504 2070 584
rect 2082 504 2086 544
rect 2090 504 2092 544
rect 2163 504 2165 544
rect 2169 540 2185 544
rect 2169 504 2171 540
rect 2183 504 2185 540
rect 2189 504 2191 544
rect 2203 504 2205 544
rect 2209 504 2211 544
rect 2268 504 2270 544
rect 2274 504 2278 544
rect 2290 504 2292 584
rect 2296 504 2300 584
rect 2304 504 2306 584
rect 2354 504 2356 584
rect 2360 504 2364 584
rect 2368 504 2370 584
rect 2382 504 2386 544
rect 2390 504 2392 544
rect 2449 504 2451 544
rect 2455 504 2457 544
rect 2469 504 2471 544
rect 2475 540 2491 544
rect 2475 504 2477 540
rect 2489 504 2491 540
rect 2495 504 2497 544
rect 2549 504 2551 544
rect 2555 504 2557 544
rect 2569 504 2571 544
rect 2575 540 2591 544
rect 2575 504 2577 540
rect 2589 504 2591 540
rect 2595 504 2597 544
rect 2663 504 2665 544
rect 2669 504 2671 544
rect 2709 504 2711 544
rect 2715 504 2717 544
rect 2729 504 2731 544
rect 2735 540 2751 544
rect 2735 504 2737 540
rect 2749 504 2751 540
rect 2755 504 2757 544
rect 2813 504 2815 584
rect 2819 544 2828 584
rect 2819 504 2821 544
rect 2833 504 2835 544
rect 2839 504 2849 544
rect 2853 504 2855 544
rect 2867 504 2869 544
rect 2873 504 2881 544
rect 2885 504 2887 544
rect 2899 504 2901 544
rect 2905 504 2907 544
rect 2945 504 2947 544
rect 2951 504 2955 544
rect 2959 524 2970 544
rect 2996 524 3005 584
rect 2959 504 2961 524
rect 2973 504 2975 524
rect 2979 504 2983 524
rect 2987 504 2991 524
rect 3003 504 3005 524
rect 3009 504 3011 584
rect 3054 504 3056 584
rect 3060 504 3064 584
rect 3068 504 3070 584
rect 3082 504 3086 544
rect 3090 504 3092 544
rect 3149 504 3151 544
rect 3155 504 3157 544
rect 3209 504 3211 544
rect 3215 504 3217 544
rect 3269 504 3271 544
rect 3275 504 3277 544
rect 3289 504 3291 544
rect 3295 540 3311 544
rect 3295 504 3297 540
rect 3309 504 3311 540
rect 3315 504 3317 544
rect 3383 504 3385 544
rect 3389 504 3391 544
rect 3443 504 3445 544
rect 3449 504 3451 544
rect 3463 504 3465 544
rect 3469 504 3471 544
rect 3528 504 3530 544
rect 3534 504 3538 544
rect 3550 504 3552 584
rect 3556 504 3560 584
rect 3564 504 3566 584
rect 3613 504 3615 584
rect 3619 544 3628 584
rect 3619 504 3621 544
rect 3633 504 3635 544
rect 3639 504 3649 544
rect 3653 504 3655 544
rect 3667 504 3669 544
rect 3673 504 3681 544
rect 3685 504 3687 544
rect 3699 504 3701 544
rect 3705 504 3707 544
rect 3745 504 3747 544
rect 3751 504 3755 544
rect 3759 524 3770 544
rect 3796 524 3805 584
rect 3759 504 3761 524
rect 3773 504 3775 524
rect 3779 504 3783 524
rect 3787 504 3791 524
rect 3803 504 3805 524
rect 3809 504 3811 584
rect 3854 504 3856 584
rect 3860 504 3864 584
rect 3868 504 3870 584
rect 3882 504 3886 544
rect 3890 504 3892 544
rect 3963 504 3965 544
rect 3969 504 3971 544
rect 3983 504 3985 544
rect 3989 504 3991 544
rect 4029 504 4031 584
rect 4035 524 4044 584
rect 4212 544 4221 584
rect 4070 524 4081 544
rect 4035 504 4037 524
rect 4049 504 4053 524
rect 4057 504 4061 524
rect 4065 504 4067 524
rect 4079 504 4081 524
rect 4085 504 4089 544
rect 4093 504 4095 544
rect 4133 504 4135 544
rect 4139 504 4141 544
rect 4153 504 4155 544
rect 4159 504 4167 544
rect 4171 504 4173 544
rect 4185 504 4187 544
rect 4191 504 4201 544
rect 4205 504 4207 544
rect 4219 504 4221 544
rect 4225 504 4227 584
rect 4269 504 4271 544
rect 4275 504 4277 544
rect 4289 504 4291 544
rect 4295 504 4297 544
rect 4349 504 4351 544
rect 4355 504 4357 544
rect 4369 504 4371 544
rect 4375 504 4377 544
rect 4448 504 4450 544
rect 4454 504 4458 544
rect 4470 504 4472 584
rect 4476 504 4480 584
rect 4484 504 4486 584
rect 4533 504 4535 584
rect 4539 544 4548 584
rect 4539 504 4541 544
rect 4553 504 4555 544
rect 4559 504 4569 544
rect 4573 504 4575 544
rect 4587 504 4589 544
rect 4593 504 4601 544
rect 4605 504 4607 544
rect 4619 504 4621 544
rect 4625 504 4627 544
rect 4665 504 4667 544
rect 4671 504 4675 544
rect 4679 524 4690 544
rect 4716 524 4725 584
rect 4679 504 4681 524
rect 4693 504 4695 524
rect 4699 504 4703 524
rect 4707 504 4711 524
rect 4723 504 4725 524
rect 4729 504 4731 584
rect 29 436 31 476
rect 35 436 37 476
rect 49 436 51 476
rect 55 436 57 476
rect 109 436 111 476
rect 115 436 117 476
rect 129 436 131 476
rect 135 436 137 476
rect 203 436 205 476
rect 209 436 211 476
rect 223 436 225 476
rect 229 436 231 476
rect 283 436 285 476
rect 289 436 291 476
rect 303 436 305 476
rect 309 436 311 476
rect 359 396 361 476
rect 365 396 367 476
rect 379 436 383 476
rect 387 436 391 476
rect 403 436 405 476
rect 409 436 411 476
rect 463 436 465 476
rect 469 436 471 476
rect 483 436 485 476
rect 489 436 491 476
rect 543 436 545 476
rect 549 440 551 476
rect 563 440 565 476
rect 549 436 565 440
rect 569 436 571 476
rect 583 436 585 476
rect 589 436 591 476
rect 643 396 645 476
rect 649 464 665 476
rect 649 396 651 464
rect 663 396 665 464
rect 669 398 671 476
rect 683 398 685 476
rect 669 396 685 398
rect 689 410 691 476
rect 703 410 705 476
rect 689 396 705 410
rect 709 398 711 476
rect 709 396 723 398
rect 775 396 777 476
rect 781 396 785 476
rect 789 396 791 476
rect 843 436 845 476
rect 849 436 851 476
rect 863 436 865 476
rect 869 436 871 476
rect 909 436 911 476
rect 915 436 917 476
rect 929 436 931 476
rect 935 436 937 476
rect 1003 436 1005 476
rect 1009 436 1011 476
rect 1023 436 1025 476
rect 1029 436 1031 476
rect 1083 436 1085 476
rect 1089 436 1091 476
rect 1103 436 1105 476
rect 1109 436 1111 476
rect 1163 396 1165 476
rect 1169 464 1185 476
rect 1169 396 1171 464
rect 1183 396 1185 464
rect 1189 398 1191 476
rect 1203 398 1205 476
rect 1189 396 1205 398
rect 1209 410 1211 476
rect 1223 410 1225 476
rect 1209 396 1225 410
rect 1229 398 1231 476
rect 1229 396 1243 398
rect 1274 396 1276 476
rect 1280 396 1284 476
rect 1288 396 1290 476
rect 1302 436 1306 476
rect 1310 436 1312 476
rect 1395 396 1397 476
rect 1401 396 1405 476
rect 1409 396 1411 476
rect 1454 396 1456 476
rect 1460 396 1464 476
rect 1468 396 1470 476
rect 1482 436 1486 476
rect 1490 436 1492 476
rect 1549 436 1551 476
rect 1555 436 1557 476
rect 1623 396 1625 476
rect 1629 396 1631 476
rect 1643 396 1645 476
rect 1649 408 1651 476
rect 1663 408 1665 476
rect 1649 396 1665 408
rect 1669 404 1671 476
rect 1709 436 1711 476
rect 1715 436 1717 476
rect 1769 436 1771 476
rect 1775 436 1777 476
rect 1789 436 1791 476
rect 1795 440 1797 476
rect 1809 440 1811 476
rect 1795 436 1811 440
rect 1815 436 1817 476
rect 1669 396 1683 404
rect 1869 404 1871 476
rect 1857 396 1871 404
rect 1875 408 1877 476
rect 1889 408 1891 476
rect 1875 396 1891 408
rect 1895 396 1897 476
rect 1909 396 1911 476
rect 1915 396 1917 476
rect 1969 436 1971 476
rect 1975 436 1977 476
rect 1989 436 1991 476
rect 1995 436 1997 476
rect 2049 436 2051 476
rect 2055 436 2057 476
rect 2069 436 2071 476
rect 2075 436 2077 476
rect 2129 436 2131 476
rect 2135 436 2137 476
rect 2149 436 2151 476
rect 2155 436 2157 476
rect 2235 396 2237 476
rect 2241 396 2245 476
rect 2249 396 2251 476
rect 2303 436 2305 476
rect 2309 436 2311 476
rect 2323 436 2325 476
rect 2329 436 2331 476
rect 2369 396 2371 476
rect 2375 396 2379 476
rect 2383 396 2385 476
rect 2449 436 2451 476
rect 2455 436 2457 476
rect 2469 436 2471 476
rect 2475 440 2477 476
rect 2489 440 2491 476
rect 2475 436 2491 440
rect 2495 436 2497 476
rect 2563 436 2565 476
rect 2569 436 2571 476
rect 2623 436 2625 476
rect 2629 440 2631 476
rect 2643 440 2645 476
rect 2629 436 2645 440
rect 2649 436 2651 476
rect 2663 436 2665 476
rect 2669 436 2671 476
rect 2709 404 2711 476
rect 2697 396 2711 404
rect 2715 408 2717 476
rect 2729 408 2731 476
rect 2715 396 2731 408
rect 2735 396 2737 476
rect 2749 396 2751 476
rect 2755 396 2757 476
rect 2809 396 2811 476
rect 2815 396 2819 476
rect 2823 396 2825 476
rect 2903 436 2905 476
rect 2909 436 2911 476
rect 2923 436 2925 476
rect 2929 436 2931 476
rect 2988 436 2990 476
rect 2994 436 2998 476
rect 3010 396 3012 476
rect 3016 396 3020 476
rect 3024 396 3026 476
rect 3088 436 3090 476
rect 3094 436 3098 476
rect 3110 396 3112 476
rect 3116 396 3120 476
rect 3124 396 3126 476
rect 3195 396 3197 476
rect 3201 396 3205 476
rect 3209 396 3211 476
rect 3263 436 3265 476
rect 3269 436 3271 476
rect 3328 436 3330 476
rect 3334 436 3338 476
rect 3350 396 3352 476
rect 3356 396 3360 476
rect 3364 396 3366 476
rect 3423 396 3425 476
rect 3429 396 3431 476
rect 3443 396 3445 476
rect 3449 408 3451 476
rect 3463 408 3465 476
rect 3449 396 3465 408
rect 3469 404 3471 476
rect 3469 396 3483 404
rect 3535 396 3537 476
rect 3541 396 3545 476
rect 3549 396 3551 476
rect 3589 396 3591 476
rect 3595 396 3601 476
rect 3605 397 3607 476
rect 3619 397 3621 476
rect 3605 396 3621 397
rect 3625 397 3627 476
rect 3689 436 3691 476
rect 3695 436 3697 476
rect 3709 436 3711 476
rect 3715 436 3717 476
rect 3769 436 3771 476
rect 3775 436 3777 476
rect 3789 436 3791 476
rect 3795 436 3797 476
rect 3868 436 3870 476
rect 3874 436 3878 476
rect 3625 396 3639 397
rect 3890 396 3892 476
rect 3896 396 3900 476
rect 3904 396 3906 476
rect 3963 436 3965 476
rect 3969 436 3971 476
rect 4023 436 4025 476
rect 4029 436 4031 476
rect 4069 396 4071 476
rect 4075 456 4077 476
rect 4089 456 4093 476
rect 4097 456 4101 476
rect 4105 456 4107 476
rect 4119 456 4121 476
rect 4075 396 4084 456
rect 4110 436 4121 456
rect 4125 436 4129 476
rect 4133 436 4135 476
rect 4173 436 4175 476
rect 4179 436 4181 476
rect 4193 436 4195 476
rect 4199 436 4207 476
rect 4211 436 4213 476
rect 4225 436 4227 476
rect 4231 436 4241 476
rect 4245 436 4247 476
rect 4259 436 4261 476
rect 4252 396 4261 436
rect 4265 396 4267 476
rect 4323 436 4325 476
rect 4329 436 4331 476
rect 4343 436 4345 476
rect 4349 436 4351 476
rect 4408 436 4410 476
rect 4414 436 4418 476
rect 4430 396 4432 476
rect 4436 396 4440 476
rect 4444 396 4446 476
rect 4503 436 4505 476
rect 4509 436 4511 476
rect 4549 396 4551 476
rect 4555 456 4557 476
rect 4569 456 4573 476
rect 4577 456 4581 476
rect 4585 456 4587 476
rect 4599 456 4601 476
rect 4555 396 4564 456
rect 4590 436 4601 456
rect 4605 436 4609 476
rect 4613 436 4615 476
rect 4653 436 4655 476
rect 4659 436 4661 476
rect 4673 436 4675 476
rect 4679 436 4687 476
rect 4691 436 4693 476
rect 4705 436 4707 476
rect 4711 436 4721 476
rect 4725 436 4727 476
rect 4739 436 4741 476
rect 4732 396 4741 436
rect 4745 396 4747 476
rect 117 96 131 104
rect 43 24 45 64
rect 49 60 65 64
rect 49 24 51 60
rect 63 24 65 60
rect 69 24 71 64
rect 83 24 85 64
rect 89 24 91 64
rect 129 24 131 96
rect 135 92 151 104
rect 135 24 137 92
rect 149 24 151 92
rect 155 24 157 104
rect 169 24 171 104
rect 175 24 177 104
rect 248 24 250 64
rect 254 24 258 64
rect 270 24 272 104
rect 276 24 280 104
rect 284 24 286 104
rect 334 24 336 104
rect 340 24 344 104
rect 348 24 350 104
rect 617 96 631 104
rect 362 24 366 64
rect 370 24 372 64
rect 443 24 445 64
rect 449 60 465 64
rect 449 24 451 60
rect 463 24 465 60
rect 469 24 471 64
rect 483 24 485 64
rect 489 24 491 64
rect 529 24 531 64
rect 535 24 537 64
rect 549 24 551 64
rect 555 60 571 64
rect 555 24 557 60
rect 569 24 571 60
rect 575 24 577 64
rect 629 24 631 96
rect 635 92 651 104
rect 635 24 637 92
rect 649 24 651 92
rect 655 24 657 104
rect 669 24 671 104
rect 675 24 677 104
rect 743 24 745 104
rect 749 24 751 104
rect 763 24 765 104
rect 769 92 785 104
rect 769 24 771 92
rect 783 24 785 92
rect 789 96 803 104
rect 789 24 791 96
rect 829 24 831 64
rect 835 24 837 64
rect 908 24 910 64
rect 914 24 918 64
rect 930 24 932 104
rect 936 24 940 104
rect 944 24 946 104
rect 1003 24 1005 64
rect 1009 24 1011 64
rect 1054 24 1056 104
rect 1060 24 1064 104
rect 1068 24 1070 104
rect 1082 24 1086 64
rect 1090 24 1092 64
rect 1154 24 1156 104
rect 1160 24 1164 104
rect 1168 24 1170 104
rect 1182 24 1186 64
rect 1190 24 1192 64
rect 1249 24 1251 64
rect 1255 24 1257 64
rect 1269 24 1271 64
rect 1275 60 1291 64
rect 1275 24 1277 60
rect 1289 24 1291 60
rect 1295 24 1297 64
rect 1349 24 1351 64
rect 1355 24 1357 64
rect 1369 24 1371 64
rect 1375 60 1391 64
rect 1375 24 1377 60
rect 1389 24 1391 60
rect 1395 24 1397 64
rect 1463 24 1465 104
rect 1469 24 1471 104
rect 1483 24 1485 104
rect 1489 92 1505 104
rect 1489 24 1491 92
rect 1503 24 1505 92
rect 1509 96 1523 104
rect 1509 24 1511 96
rect 1549 24 1551 64
rect 1555 24 1557 64
rect 1569 24 1571 64
rect 1575 60 1591 64
rect 1575 24 1577 60
rect 1589 24 1591 60
rect 1595 24 1597 64
rect 1663 24 1665 104
rect 1669 24 1671 104
rect 1683 24 1685 104
rect 1689 92 1705 104
rect 1689 24 1691 92
rect 1703 24 1705 92
rect 1709 96 1723 104
rect 1709 24 1711 96
rect 1749 24 1751 64
rect 1755 24 1757 64
rect 1769 24 1771 64
rect 1775 60 1791 64
rect 1775 24 1777 60
rect 1789 24 1791 60
rect 1795 24 1797 64
rect 1849 24 1851 64
rect 1855 24 1857 64
rect 1869 24 1871 64
rect 1875 24 1877 64
rect 1929 24 1931 64
rect 1935 24 1939 64
rect 1951 24 1953 104
rect 1957 24 1959 104
rect 2019 24 2021 104
rect 2025 24 2027 104
rect 2039 24 2043 64
rect 2047 24 2051 64
rect 2063 24 2065 64
rect 2069 24 2071 64
rect 2109 24 2111 64
rect 2115 24 2119 64
rect 2131 24 2133 104
rect 2137 24 2139 104
rect 2277 102 2291 104
rect 2189 24 2191 64
rect 2195 24 2197 64
rect 2209 24 2211 64
rect 2215 60 2231 64
rect 2215 24 2217 60
rect 2229 24 2231 60
rect 2235 24 2237 64
rect 2289 24 2291 102
rect 2295 90 2311 104
rect 2295 24 2297 90
rect 2309 24 2311 90
rect 2315 102 2331 104
rect 2315 24 2317 102
rect 2329 24 2331 102
rect 2335 36 2337 104
rect 2349 36 2351 104
rect 2335 24 2351 36
rect 2355 24 2357 104
rect 2414 24 2416 104
rect 2420 24 2424 104
rect 2428 24 2430 104
rect 2442 24 2446 64
rect 2450 24 2452 64
rect 2523 24 2525 104
rect 2529 24 2531 104
rect 2543 24 2545 104
rect 2549 92 2565 104
rect 2549 24 2551 92
rect 2563 24 2565 92
rect 2569 96 2583 104
rect 2569 24 2571 96
rect 2614 24 2616 104
rect 2620 24 2624 104
rect 2628 24 2630 104
rect 2642 24 2646 64
rect 2650 24 2652 64
rect 2709 24 2711 64
rect 2715 24 2717 64
rect 2769 24 2771 64
rect 2775 24 2777 64
rect 2789 24 2791 64
rect 2795 60 2811 64
rect 2795 24 2797 60
rect 2809 24 2811 60
rect 2815 24 2817 64
rect 2869 24 2871 64
rect 2875 24 2877 64
rect 2933 24 2935 104
rect 2939 64 2948 104
rect 2939 24 2941 64
rect 2953 24 2955 64
rect 2959 24 2969 64
rect 2973 24 2975 64
rect 2987 24 2989 64
rect 2993 24 3001 64
rect 3005 24 3007 64
rect 3019 24 3021 64
rect 3025 24 3027 64
rect 3065 24 3067 64
rect 3071 24 3075 64
rect 3079 44 3090 64
rect 3116 44 3125 104
rect 3079 24 3081 44
rect 3093 24 3095 44
rect 3099 24 3103 44
rect 3107 24 3111 44
rect 3123 24 3125 44
rect 3129 24 3131 104
rect 3169 24 3171 64
rect 3175 24 3177 64
rect 3243 24 3245 64
rect 3249 24 3251 64
rect 3293 24 3295 104
rect 3299 64 3308 104
rect 3299 24 3301 64
rect 3313 24 3315 64
rect 3319 24 3329 64
rect 3333 24 3335 64
rect 3347 24 3349 64
rect 3353 24 3361 64
rect 3365 24 3367 64
rect 3379 24 3381 64
rect 3385 24 3387 64
rect 3425 24 3427 64
rect 3431 24 3435 64
rect 3439 44 3450 64
rect 3476 44 3485 104
rect 3439 24 3441 44
rect 3453 24 3455 44
rect 3459 24 3463 44
rect 3467 24 3471 44
rect 3483 24 3485 44
rect 3489 24 3491 104
rect 3555 24 3557 104
rect 3561 24 3565 104
rect 3569 24 3571 104
rect 3609 24 3611 104
rect 3615 44 3624 104
rect 3792 64 3801 104
rect 3650 44 3661 64
rect 3615 24 3617 44
rect 3629 24 3633 44
rect 3637 24 3641 44
rect 3645 24 3647 44
rect 3659 24 3661 44
rect 3665 24 3669 64
rect 3673 24 3675 64
rect 3713 24 3715 64
rect 3719 24 3721 64
rect 3733 24 3735 64
rect 3739 24 3747 64
rect 3751 24 3753 64
rect 3765 24 3767 64
rect 3771 24 3781 64
rect 3785 24 3787 64
rect 3799 24 3801 64
rect 3805 24 3807 104
rect 3849 24 3851 64
rect 3855 24 3857 64
rect 3914 24 3916 104
rect 3920 24 3924 104
rect 3928 24 3930 104
rect 3942 24 3946 64
rect 3950 24 3952 64
rect 4009 24 4011 104
rect 4015 24 4019 104
rect 4023 24 4025 104
rect 4089 24 4091 104
rect 4095 24 4099 104
rect 4103 24 4105 104
rect 4195 24 4197 104
rect 4201 24 4205 104
rect 4209 24 4211 104
rect 4254 24 4256 104
rect 4260 24 4264 104
rect 4268 24 4270 104
rect 4282 24 4286 64
rect 4290 24 4292 64
rect 4363 24 4365 64
rect 4369 24 4371 64
rect 4383 24 4385 64
rect 4389 24 4391 64
rect 4443 24 4445 64
rect 4449 24 4451 64
rect 4489 24 4491 104
rect 4495 24 4499 104
rect 4503 24 4505 104
rect 4569 24 4571 64
rect 4575 24 4577 64
rect 4589 24 4591 64
rect 4595 24 4597 64
rect 4663 24 4665 64
rect 4669 24 4671 64
rect 4709 24 4711 64
rect 4715 24 4717 64
rect 4729 24 4731 64
rect 4735 24 4737 64
<< ndcontact >>
rect 38 4536 50 4556
rect 60 4516 72 4556
rect 88 4516 100 4556
rect 154 4498 166 4556
rect 190 4496 202 4556
rect 218 4496 230 4556
rect 254 4498 266 4556
rect 354 4498 366 4556
rect 390 4496 402 4556
rect 420 4516 432 4556
rect 448 4516 460 4556
rect 470 4536 482 4556
rect 517 4516 529 4556
rect 537 4528 549 4556
rect 557 4516 569 4556
rect 577 4516 589 4556
rect 617 4516 629 4556
rect 637 4528 649 4556
rect 657 4516 669 4556
rect 677 4516 689 4556
rect 754 4498 766 4556
rect 790 4496 802 4556
rect 818 4496 830 4556
rect 854 4498 866 4556
rect 919 4516 931 4556
rect 949 4516 961 4556
rect 998 4496 1010 4556
rect 1034 4498 1046 4556
rect 1100 4516 1112 4556
rect 1128 4516 1140 4556
rect 1150 4536 1162 4556
rect 1219 4516 1231 4556
rect 1249 4516 1261 4556
rect 1291 4536 1303 4556
rect 1311 4536 1323 4556
rect 1331 4536 1343 4556
rect 1371 4516 1383 4556
rect 1391 4516 1403 4556
rect 1411 4528 1423 4556
rect 1431 4516 1443 4556
rect 1479 4516 1491 4556
rect 1509 4516 1521 4556
rect 1537 4536 1549 4556
rect 1557 4536 1569 4556
rect 1577 4536 1589 4556
rect 1618 4496 1630 4556
rect 1654 4498 1666 4556
rect 1738 4536 1750 4556
rect 1760 4516 1772 4556
rect 1788 4516 1800 4556
rect 1817 4536 1829 4556
rect 1837 4536 1849 4556
rect 1891 4536 1903 4556
rect 1911 4536 1923 4556
rect 1940 4516 1952 4556
rect 1968 4516 1980 4556
rect 1990 4536 2002 4556
rect 2037 4536 2049 4556
rect 2057 4536 2069 4556
rect 2077 4536 2089 4556
rect 2117 4536 2129 4556
rect 2137 4536 2149 4556
rect 2177 4516 2189 4556
rect 2197 4528 2209 4556
rect 2217 4516 2229 4556
rect 2237 4516 2249 4556
rect 2291 4516 2303 4556
rect 2311 4516 2323 4544
rect 2331 4516 2343 4556
rect 2351 4526 2363 4556
rect 2371 4516 2383 4556
rect 2397 4536 2409 4556
rect 2417 4536 2429 4556
rect 2437 4536 2449 4556
rect 2457 4516 2469 4556
rect 2500 4516 2512 4556
rect 2528 4516 2540 4556
rect 2550 4536 2562 4556
rect 2632 4516 2644 4556
rect 2660 4516 2672 4556
rect 2688 4516 2700 4556
rect 2721 4516 2733 4556
rect 2741 4536 2753 4556
rect 2773 4536 2785 4556
rect 2803 4536 2815 4556
rect 2825 4536 2837 4556
rect 2851 4536 2863 4556
rect 2879 4536 2891 4556
rect 2909 4536 2921 4556
rect 2931 4516 2943 4556
rect 2971 4536 2983 4556
rect 2991 4536 3003 4556
rect 3031 4516 3043 4556
rect 3051 4516 3063 4556
rect 3071 4528 3083 4556
rect 3091 4516 3103 4556
rect 3131 4536 3143 4556
rect 3151 4536 3163 4556
rect 3171 4536 3183 4556
rect 3211 4516 3223 4556
rect 3231 4516 3243 4556
rect 3251 4528 3263 4556
rect 3271 4516 3283 4556
rect 3311 4536 3323 4556
rect 3331 4536 3343 4556
rect 3351 4536 3363 4556
rect 3391 4536 3403 4556
rect 3411 4536 3423 4556
rect 3437 4516 3449 4556
rect 3459 4536 3471 4556
rect 3489 4536 3501 4556
rect 3517 4536 3529 4556
rect 3543 4536 3555 4556
rect 3565 4536 3577 4556
rect 3595 4536 3607 4556
rect 3627 4536 3639 4556
rect 3647 4516 3659 4556
rect 3677 4516 3689 4556
rect 3697 4528 3709 4556
rect 3717 4516 3729 4556
rect 3737 4516 3749 4556
rect 3779 4516 3791 4556
rect 3809 4516 3821 4556
rect 3871 4516 3883 4556
rect 3891 4516 3903 4556
rect 3911 4516 3923 4556
rect 3931 4516 3943 4556
rect 3951 4516 3963 4556
rect 3971 4516 3983 4556
rect 3991 4516 4003 4556
rect 4011 4516 4023 4556
rect 4031 4516 4043 4556
rect 4069 4516 4081 4556
rect 4089 4516 4101 4556
rect 4111 4536 4123 4556
rect 4139 4516 4151 4556
rect 4169 4516 4181 4556
rect 4217 4536 4229 4556
rect 4237 4536 4249 4556
rect 4277 4516 4289 4556
rect 4297 4528 4309 4556
rect 4317 4516 4329 4556
rect 4337 4516 4349 4556
rect 4377 4516 4389 4556
rect 4399 4536 4411 4556
rect 4429 4536 4441 4556
rect 4457 4536 4469 4556
rect 4483 4536 4495 4556
rect 4505 4536 4517 4556
rect 4535 4536 4547 4556
rect 4567 4536 4579 4556
rect 4587 4516 4599 4556
rect 4617 4536 4629 4556
rect 4639 4516 4651 4556
rect 4659 4516 4671 4556
rect 4699 4516 4711 4556
rect 4729 4516 4741 4556
rect 39 4104 51 4144
rect 69 4104 81 4144
rect 100 4104 112 4144
rect 128 4104 140 4144
rect 150 4104 162 4124
rect 219 4104 231 4144
rect 249 4104 261 4144
rect 291 4104 303 4124
rect 311 4104 323 4124
rect 331 4104 343 4124
rect 371 4104 383 4144
rect 391 4104 403 4144
rect 411 4104 423 4132
rect 431 4104 443 4144
rect 457 4104 469 4144
rect 477 4104 489 4132
rect 497 4104 509 4144
rect 517 4104 529 4144
rect 571 4104 583 4124
rect 591 4104 603 4124
rect 638 4104 650 4124
rect 660 4104 672 4144
rect 688 4104 700 4144
rect 731 4104 743 4124
rect 751 4104 763 4124
rect 778 4104 790 4164
rect 814 4104 826 4162
rect 912 4104 924 4144
rect 940 4104 952 4144
rect 968 4104 980 4144
rect 1034 4104 1046 4162
rect 1070 4104 1082 4164
rect 1098 4104 1110 4164
rect 1134 4104 1146 4162
rect 1219 4104 1231 4144
rect 1249 4104 1261 4144
rect 1314 4104 1326 4162
rect 1350 4104 1362 4164
rect 1399 4104 1411 4144
rect 1429 4104 1441 4144
rect 1458 4104 1470 4164
rect 1494 4104 1506 4162
rect 1571 4104 1583 4124
rect 1591 4104 1603 4124
rect 1611 4104 1623 4124
rect 1651 4104 1663 4124
rect 1671 4104 1683 4124
rect 1691 4104 1703 4124
rect 1717 4104 1729 4144
rect 1737 4104 1749 4132
rect 1757 4104 1769 4144
rect 1777 4104 1789 4144
rect 1839 4104 1851 4144
rect 1869 4104 1881 4144
rect 1897 4104 1909 4124
rect 1917 4104 1929 4124
rect 1958 4104 1970 4164
rect 1994 4104 2006 4162
rect 2058 4104 2070 4164
rect 2094 4104 2106 4162
rect 2161 4104 2173 4144
rect 2181 4104 2193 4124
rect 2213 4104 2225 4124
rect 2243 4104 2255 4124
rect 2265 4104 2277 4124
rect 2291 4104 2303 4124
rect 2319 4104 2331 4124
rect 2349 4104 2361 4124
rect 2371 4104 2383 4144
rect 2397 4104 2409 4124
rect 2419 4104 2431 4144
rect 2439 4104 2451 4144
rect 2491 4104 2503 4124
rect 2511 4104 2523 4124
rect 2551 4104 2563 4124
rect 2571 4104 2583 4124
rect 2591 4104 2603 4124
rect 2617 4104 2629 4144
rect 2639 4104 2651 4124
rect 2669 4104 2681 4124
rect 2697 4104 2709 4124
rect 2723 4104 2735 4124
rect 2745 4104 2757 4124
rect 2775 4104 2787 4124
rect 2807 4104 2819 4124
rect 2827 4104 2839 4144
rect 2857 4104 2869 4124
rect 2877 4104 2889 4124
rect 2931 4104 2943 4124
rect 2951 4104 2963 4124
rect 2971 4104 2983 4124
rect 2997 4104 3009 4144
rect 3017 4104 3029 4132
rect 3037 4104 3049 4144
rect 3057 4104 3069 4144
rect 3099 4104 3111 4144
rect 3129 4104 3141 4144
rect 3199 4104 3211 4144
rect 3229 4104 3241 4144
rect 3279 4104 3291 4144
rect 3309 4104 3321 4144
rect 3337 4104 3349 4124
rect 3357 4104 3369 4124
rect 3377 4104 3389 4124
rect 3421 4104 3433 4144
rect 3441 4104 3453 4124
rect 3473 4104 3485 4124
rect 3503 4104 3515 4124
rect 3525 4104 3537 4124
rect 3551 4104 3563 4124
rect 3579 4104 3591 4124
rect 3609 4104 3621 4124
rect 3631 4104 3643 4144
rect 3679 4104 3691 4144
rect 3709 4104 3721 4144
rect 3737 4104 3749 4124
rect 3757 4104 3769 4124
rect 3777 4104 3789 4124
rect 3817 4104 3829 4144
rect 3839 4104 3851 4124
rect 3869 4104 3881 4124
rect 3897 4104 3909 4124
rect 3923 4104 3935 4124
rect 3945 4104 3957 4124
rect 3975 4104 3987 4124
rect 4007 4104 4019 4124
rect 4027 4104 4039 4144
rect 4057 4104 4069 4124
rect 4077 4104 4089 4124
rect 4097 4104 4109 4124
rect 4158 4104 4170 4124
rect 4180 4104 4192 4144
rect 4208 4104 4220 4144
rect 4237 4104 4249 4124
rect 4259 4104 4271 4144
rect 4279 4104 4291 4144
rect 4331 4104 4343 4124
rect 4351 4104 4363 4124
rect 4371 4104 4383 4124
rect 4418 4104 4430 4124
rect 4440 4104 4452 4144
rect 4468 4104 4480 4144
rect 4497 4104 4509 4144
rect 4519 4104 4531 4124
rect 4549 4104 4561 4124
rect 4577 4104 4589 4124
rect 4603 4104 4615 4124
rect 4625 4104 4637 4124
rect 4655 4104 4667 4124
rect 4687 4104 4699 4124
rect 4707 4104 4719 4144
rect 39 4036 51 4076
rect 69 4036 81 4076
rect 99 4036 111 4076
rect 129 4036 141 4076
rect 199 4036 211 4076
rect 229 4036 241 4076
rect 271 4036 283 4076
rect 291 4036 303 4076
rect 311 4048 323 4076
rect 331 4036 343 4076
rect 360 4036 372 4076
rect 388 4036 400 4076
rect 410 4056 422 4076
rect 471 4056 483 4076
rect 491 4056 503 4076
rect 511 4056 523 4076
rect 539 4036 551 4076
rect 569 4036 581 4076
rect 617 4036 629 4076
rect 637 4048 649 4076
rect 657 4036 669 4076
rect 677 4036 689 4076
rect 754 4018 766 4076
rect 790 4016 802 4076
rect 818 4016 830 4076
rect 854 4018 866 4076
rect 931 4036 943 4076
rect 951 4036 963 4076
rect 971 4048 983 4076
rect 991 4036 1003 4076
rect 1017 4036 1029 4076
rect 1037 4048 1049 4076
rect 1057 4036 1069 4076
rect 1077 4036 1089 4076
rect 1131 4056 1143 4076
rect 1151 4056 1163 4076
rect 1214 4018 1226 4076
rect 1250 4016 1262 4076
rect 1277 4056 1289 4076
rect 1297 4056 1309 4076
rect 1338 4016 1350 4076
rect 1374 4018 1386 4076
rect 1438 4016 1450 4076
rect 1474 4018 1486 4076
rect 1539 4036 1551 4076
rect 1569 4036 1581 4076
rect 1631 4056 1643 4076
rect 1651 4056 1663 4076
rect 1671 4056 1683 4076
rect 1721 4036 1733 4076
rect 1741 4036 1753 4076
rect 1771 4036 1783 4076
rect 1811 4036 1823 4076
rect 1831 4036 1843 4076
rect 1851 4048 1863 4076
rect 1871 4036 1883 4076
rect 1897 4056 1909 4076
rect 1917 4056 1929 4076
rect 1937 4056 1949 4076
rect 1991 4056 2003 4076
rect 2011 4056 2023 4076
rect 2037 4036 2049 4076
rect 2057 4048 2069 4076
rect 2077 4036 2089 4076
rect 2097 4036 2109 4076
rect 2137 4056 2149 4076
rect 2157 4056 2169 4076
rect 2199 4036 2211 4076
rect 2229 4036 2241 4076
rect 2278 4016 2290 4076
rect 2314 4018 2326 4076
rect 2377 4056 2389 4076
rect 2399 4036 2411 4076
rect 2419 4036 2431 4076
rect 2457 4036 2469 4076
rect 2477 4036 2489 4076
rect 2497 4036 2509 4076
rect 2517 4036 2529 4076
rect 2537 4036 2549 4076
rect 2557 4036 2569 4076
rect 2577 4036 2589 4076
rect 2597 4036 2609 4076
rect 2617 4036 2629 4076
rect 2661 4036 2673 4076
rect 2681 4056 2693 4076
rect 2713 4056 2725 4076
rect 2743 4056 2755 4076
rect 2765 4056 2777 4076
rect 2791 4056 2803 4076
rect 2819 4056 2831 4076
rect 2849 4056 2861 4076
rect 2871 4036 2883 4076
rect 2897 4056 2909 4076
rect 2917 4056 2929 4076
rect 2957 4036 2969 4076
rect 2977 4048 2989 4076
rect 2997 4036 3009 4076
rect 3017 4036 3029 4076
rect 3057 4056 3069 4076
rect 3077 4056 3089 4076
rect 3097 4056 3109 4076
rect 3139 4036 3151 4076
rect 3169 4036 3181 4076
rect 3238 4056 3250 4076
rect 3260 4036 3272 4076
rect 3288 4036 3300 4076
rect 3317 4036 3329 4076
rect 3347 4036 3359 4076
rect 3367 4036 3379 4076
rect 3431 4056 3443 4076
rect 3451 4056 3463 4076
rect 3471 4056 3483 4076
rect 3511 4056 3523 4076
rect 3531 4056 3543 4076
rect 3557 4036 3569 4076
rect 3579 4056 3591 4076
rect 3609 4056 3621 4076
rect 3637 4056 3649 4076
rect 3663 4056 3675 4076
rect 3685 4056 3697 4076
rect 3715 4056 3727 4076
rect 3747 4056 3759 4076
rect 3767 4036 3779 4076
rect 3818 4056 3830 4076
rect 3840 4036 3852 4076
rect 3868 4036 3880 4076
rect 3897 4056 3909 4076
rect 3917 4056 3929 4076
rect 3937 4056 3949 4076
rect 3991 4056 4003 4076
rect 4011 4056 4023 4076
rect 4031 4056 4043 4076
rect 4057 4036 4069 4076
rect 4087 4036 4099 4076
rect 4107 4036 4119 4076
rect 4157 4036 4169 4076
rect 4177 4048 4189 4076
rect 4197 4036 4209 4076
rect 4217 4036 4229 4076
rect 4271 4036 4283 4076
rect 4291 4036 4303 4076
rect 4311 4048 4323 4076
rect 4331 4036 4343 4076
rect 4371 4056 4383 4076
rect 4391 4056 4403 4076
rect 4417 4036 4429 4076
rect 4439 4056 4451 4076
rect 4469 4056 4481 4076
rect 4497 4056 4509 4076
rect 4523 4056 4535 4076
rect 4545 4056 4557 4076
rect 4575 4056 4587 4076
rect 4607 4056 4619 4076
rect 4627 4036 4639 4076
rect 4657 4056 4669 4076
rect 4677 4056 4689 4076
rect 31 3624 43 3644
rect 51 3624 63 3644
rect 71 3624 83 3644
rect 97 3624 109 3664
rect 117 3624 129 3652
rect 137 3624 149 3664
rect 157 3624 169 3664
rect 211 3624 223 3644
rect 231 3624 243 3644
rect 278 3624 290 3644
rect 300 3624 312 3664
rect 328 3624 340 3664
rect 381 3624 393 3664
rect 401 3624 413 3664
rect 431 3624 443 3664
rect 479 3624 491 3664
rect 509 3624 521 3664
rect 559 3624 571 3664
rect 589 3624 601 3664
rect 617 3624 629 3644
rect 637 3624 649 3644
rect 677 3624 689 3664
rect 697 3624 709 3652
rect 717 3624 729 3664
rect 737 3624 749 3664
rect 779 3624 791 3664
rect 809 3624 821 3664
rect 894 3624 906 3682
rect 930 3624 942 3684
rect 960 3624 972 3664
rect 988 3624 1000 3664
rect 1010 3624 1022 3644
rect 1058 3624 1070 3684
rect 1094 3624 1106 3682
rect 1160 3624 1172 3664
rect 1188 3624 1200 3664
rect 1210 3624 1222 3644
rect 1257 3624 1269 3644
rect 1277 3624 1289 3644
rect 1354 3624 1366 3682
rect 1390 3624 1402 3684
rect 1431 3624 1443 3644
rect 1451 3624 1463 3644
rect 1491 3624 1503 3664
rect 1511 3624 1523 3664
rect 1531 3624 1543 3652
rect 1551 3624 1563 3664
rect 1591 3624 1603 3644
rect 1611 3624 1623 3644
rect 1640 3624 1652 3664
rect 1668 3624 1680 3664
rect 1690 3624 1702 3644
rect 1737 3624 1749 3644
rect 1757 3624 1769 3644
rect 1777 3624 1789 3644
rect 1838 3624 1850 3644
rect 1860 3624 1872 3664
rect 1888 3624 1900 3664
rect 1939 3624 1951 3664
rect 1969 3624 1981 3664
rect 1997 3624 2009 3644
rect 2017 3624 2029 3644
rect 2037 3624 2049 3644
rect 2057 3624 2069 3664
rect 2097 3624 2109 3644
rect 2119 3624 2131 3664
rect 2139 3624 2151 3664
rect 2191 3624 2203 3664
rect 2211 3624 2223 3664
rect 2231 3624 2243 3664
rect 2251 3624 2263 3664
rect 2271 3624 2283 3664
rect 2291 3624 2303 3664
rect 2311 3624 2323 3664
rect 2331 3624 2343 3664
rect 2351 3624 2363 3664
rect 2381 3624 2393 3664
rect 2401 3624 2413 3644
rect 2433 3624 2445 3644
rect 2463 3624 2475 3644
rect 2485 3624 2497 3644
rect 2511 3624 2523 3644
rect 2539 3624 2551 3644
rect 2569 3624 2581 3644
rect 2591 3624 2603 3664
rect 2631 3624 2643 3664
rect 2651 3624 2663 3664
rect 2671 3624 2683 3652
rect 2691 3624 2703 3664
rect 2731 3624 2743 3644
rect 2751 3624 2763 3644
rect 2791 3624 2803 3644
rect 2811 3624 2823 3644
rect 2831 3624 2843 3644
rect 2871 3624 2883 3644
rect 2891 3624 2903 3644
rect 2911 3624 2923 3644
rect 2951 3624 2963 3644
rect 2971 3624 2983 3644
rect 2991 3624 3003 3644
rect 3017 3624 3029 3644
rect 3037 3624 3049 3644
rect 3091 3624 3103 3644
rect 3111 3624 3123 3644
rect 3137 3624 3149 3664
rect 3157 3624 3169 3652
rect 3177 3624 3189 3664
rect 3197 3624 3209 3664
rect 3258 3624 3270 3644
rect 3280 3624 3292 3664
rect 3308 3624 3320 3664
rect 3340 3624 3352 3664
rect 3368 3624 3380 3664
rect 3390 3624 3402 3644
rect 3437 3624 3449 3644
rect 3457 3624 3469 3644
rect 3497 3624 3509 3664
rect 3527 3624 3539 3664
rect 3547 3624 3559 3664
rect 3597 3624 3609 3664
rect 3617 3624 3629 3652
rect 3637 3624 3649 3664
rect 3657 3624 3669 3664
rect 3697 3624 3709 3664
rect 3717 3624 3729 3652
rect 3737 3624 3749 3664
rect 3757 3624 3769 3664
rect 3801 3624 3813 3664
rect 3821 3624 3833 3644
rect 3853 3624 3865 3644
rect 3883 3624 3895 3644
rect 3905 3624 3917 3644
rect 3931 3624 3943 3644
rect 3959 3624 3971 3644
rect 3989 3624 4001 3644
rect 4011 3624 4023 3664
rect 4037 3624 4049 3644
rect 4059 3624 4071 3664
rect 4079 3624 4091 3664
rect 4131 3624 4143 3644
rect 4151 3624 4163 3644
rect 4171 3624 4183 3644
rect 4200 3624 4212 3664
rect 4228 3624 4240 3664
rect 4250 3624 4262 3644
rect 4297 3624 4309 3664
rect 4319 3624 4331 3644
rect 4349 3624 4361 3644
rect 4377 3624 4389 3644
rect 4403 3624 4415 3644
rect 4425 3624 4437 3644
rect 4455 3624 4467 3644
rect 4487 3624 4499 3644
rect 4507 3624 4519 3664
rect 4537 3624 4549 3644
rect 4559 3624 4571 3664
rect 4579 3624 4591 3664
rect 4631 3624 4643 3644
rect 4651 3624 4663 3644
rect 4677 3624 4689 3644
rect 4697 3624 4709 3644
rect 39 3556 51 3596
rect 69 3556 81 3596
rect 101 3556 113 3596
rect 121 3576 133 3596
rect 153 3576 165 3596
rect 183 3576 195 3596
rect 205 3576 217 3596
rect 231 3576 243 3596
rect 259 3576 271 3596
rect 289 3576 301 3596
rect 311 3556 323 3596
rect 351 3576 363 3596
rect 371 3576 383 3596
rect 419 3556 431 3596
rect 449 3556 461 3596
rect 491 3556 503 3596
rect 511 3556 523 3596
rect 531 3568 543 3596
rect 551 3556 563 3596
rect 591 3556 603 3596
rect 611 3556 623 3596
rect 631 3568 643 3596
rect 651 3556 663 3596
rect 679 3556 691 3596
rect 709 3556 721 3596
rect 757 3556 769 3596
rect 777 3566 789 3596
rect 797 3556 809 3596
rect 817 3556 829 3584
rect 837 3556 849 3596
rect 877 3576 889 3596
rect 897 3576 909 3596
rect 974 3538 986 3596
rect 1010 3536 1022 3596
rect 1040 3556 1052 3596
rect 1068 3556 1080 3596
rect 1090 3576 1102 3596
rect 1137 3576 1149 3596
rect 1157 3576 1169 3596
rect 1177 3576 1189 3596
rect 1219 3556 1231 3596
rect 1249 3556 1261 3596
rect 1299 3556 1311 3596
rect 1329 3556 1341 3596
rect 1377 3556 1389 3596
rect 1397 3568 1409 3596
rect 1417 3556 1429 3596
rect 1437 3556 1449 3596
rect 1481 3556 1493 3596
rect 1501 3576 1513 3596
rect 1533 3576 1545 3596
rect 1563 3576 1575 3596
rect 1585 3576 1597 3596
rect 1611 3576 1623 3596
rect 1639 3576 1651 3596
rect 1669 3576 1681 3596
rect 1691 3556 1703 3596
rect 1739 3556 1751 3596
rect 1769 3556 1781 3596
rect 1797 3556 1809 3596
rect 1817 3568 1829 3596
rect 1837 3556 1849 3596
rect 1857 3556 1869 3596
rect 1897 3556 1909 3596
rect 1917 3556 1929 3596
rect 1979 3556 1991 3596
rect 2009 3556 2021 3596
rect 2061 3556 2073 3596
rect 2081 3556 2093 3596
rect 2111 3556 2123 3596
rect 2139 3556 2151 3596
rect 2169 3556 2181 3596
rect 2218 3536 2230 3596
rect 2254 3538 2266 3596
rect 2317 3576 2329 3596
rect 2337 3576 2349 3596
rect 2377 3576 2389 3596
rect 2397 3576 2409 3596
rect 2437 3556 2449 3596
rect 2459 3576 2471 3596
rect 2489 3576 2501 3596
rect 2517 3576 2529 3596
rect 2543 3576 2555 3596
rect 2565 3576 2577 3596
rect 2595 3576 2607 3596
rect 2627 3576 2639 3596
rect 2647 3556 2659 3596
rect 2677 3556 2689 3596
rect 2697 3568 2709 3596
rect 2717 3556 2729 3596
rect 2737 3556 2749 3596
rect 2777 3576 2789 3596
rect 2799 3556 2811 3596
rect 2819 3556 2831 3596
rect 2859 3556 2871 3596
rect 2889 3556 2901 3596
rect 2937 3556 2949 3596
rect 2959 3576 2971 3596
rect 2989 3576 3001 3596
rect 3017 3576 3029 3596
rect 3043 3576 3055 3596
rect 3065 3576 3077 3596
rect 3095 3576 3107 3596
rect 3127 3576 3139 3596
rect 3147 3556 3159 3596
rect 3191 3556 3203 3596
rect 3211 3556 3223 3596
rect 3231 3568 3243 3596
rect 3251 3556 3263 3596
rect 3291 3576 3303 3596
rect 3311 3576 3323 3596
rect 3337 3576 3349 3596
rect 3357 3576 3369 3596
rect 3377 3576 3389 3596
rect 3417 3576 3429 3596
rect 3437 3576 3449 3596
rect 3491 3576 3503 3596
rect 3511 3576 3523 3596
rect 3531 3576 3543 3596
rect 3560 3556 3572 3596
rect 3588 3556 3600 3596
rect 3610 3576 3622 3596
rect 3657 3576 3669 3596
rect 3677 3576 3689 3596
rect 3697 3576 3709 3596
rect 3717 3556 3729 3596
rect 3792 3556 3804 3596
rect 3820 3556 3832 3596
rect 3848 3556 3860 3596
rect 3899 3556 3911 3596
rect 3929 3556 3941 3596
rect 3957 3556 3969 3596
rect 3979 3576 3991 3596
rect 4009 3576 4021 3596
rect 4037 3576 4049 3596
rect 4063 3576 4075 3596
rect 4085 3576 4097 3596
rect 4115 3576 4127 3596
rect 4147 3576 4159 3596
rect 4167 3556 4179 3596
rect 4197 3556 4209 3596
rect 4219 3576 4231 3596
rect 4249 3576 4261 3596
rect 4277 3576 4289 3596
rect 4303 3576 4315 3596
rect 4325 3576 4337 3596
rect 4355 3576 4367 3596
rect 4387 3576 4399 3596
rect 4407 3556 4419 3596
rect 4451 3556 4463 3596
rect 4471 3556 4483 3596
rect 4491 3556 4503 3596
rect 4511 3556 4523 3596
rect 4531 3556 4543 3596
rect 4551 3556 4563 3596
rect 4571 3556 4583 3596
rect 4591 3556 4603 3596
rect 4611 3556 4623 3596
rect 4637 3556 4649 3596
rect 4657 3568 4669 3596
rect 4677 3556 4689 3596
rect 4697 3556 4709 3596
rect 21 3144 33 3184
rect 41 3144 53 3164
rect 73 3144 85 3164
rect 103 3144 115 3164
rect 125 3144 137 3164
rect 151 3144 163 3164
rect 179 3144 191 3164
rect 209 3144 221 3164
rect 231 3144 243 3184
rect 292 3144 304 3184
rect 320 3144 332 3184
rect 348 3144 360 3184
rect 399 3144 411 3184
rect 429 3144 441 3184
rect 457 3144 469 3184
rect 479 3144 491 3164
rect 509 3144 521 3164
rect 537 3144 549 3164
rect 563 3144 575 3164
rect 585 3144 597 3164
rect 615 3144 627 3164
rect 647 3144 659 3164
rect 667 3144 679 3184
rect 711 3144 723 3184
rect 731 3144 743 3184
rect 751 3144 763 3172
rect 771 3144 783 3184
rect 832 3144 844 3184
rect 860 3144 872 3184
rect 888 3144 900 3184
rect 919 3144 931 3184
rect 949 3144 961 3184
rect 1034 3144 1046 3202
rect 1070 3144 1082 3204
rect 1121 3144 1133 3184
rect 1141 3144 1153 3184
rect 1171 3144 1183 3184
rect 1198 3144 1210 3204
rect 1234 3144 1246 3202
rect 1297 3144 1309 3184
rect 1317 3144 1329 3172
rect 1337 3144 1349 3184
rect 1357 3144 1369 3184
rect 1399 3144 1411 3184
rect 1429 3144 1441 3184
rect 1491 3144 1503 3184
rect 1511 3144 1523 3164
rect 1531 3144 1543 3164
rect 1551 3144 1563 3164
rect 1599 3144 1611 3184
rect 1629 3144 1641 3184
rect 1657 3144 1669 3184
rect 1677 3144 1689 3172
rect 1697 3144 1709 3184
rect 1717 3144 1729 3184
rect 1771 3144 1783 3184
rect 1791 3144 1803 3184
rect 1811 3144 1823 3172
rect 1831 3144 1843 3184
rect 1859 3144 1871 3184
rect 1889 3144 1901 3184
rect 1937 3144 1949 3184
rect 1957 3144 1969 3172
rect 1977 3144 1989 3184
rect 1997 3144 2009 3184
rect 2051 3144 2063 3184
rect 2071 3144 2083 3184
rect 2091 3144 2103 3172
rect 2111 3144 2123 3184
rect 2137 3144 2149 3164
rect 2157 3144 2169 3164
rect 2197 3144 2209 3184
rect 2217 3144 2229 3172
rect 2237 3144 2249 3184
rect 2257 3144 2269 3184
rect 2311 3144 2323 3164
rect 2331 3144 2343 3164
rect 2359 3144 2371 3184
rect 2389 3144 2401 3184
rect 2437 3144 2449 3184
rect 2459 3144 2471 3164
rect 2489 3144 2501 3164
rect 2517 3144 2529 3164
rect 2543 3144 2555 3164
rect 2565 3144 2577 3164
rect 2595 3144 2607 3164
rect 2627 3144 2639 3164
rect 2647 3144 2659 3184
rect 2677 3144 2689 3164
rect 2699 3144 2711 3184
rect 2719 3144 2731 3184
rect 2757 3144 2769 3184
rect 2779 3144 2791 3164
rect 2809 3144 2821 3164
rect 2837 3144 2849 3164
rect 2863 3144 2875 3164
rect 2885 3144 2897 3164
rect 2915 3144 2927 3164
rect 2947 3144 2959 3164
rect 2967 3144 2979 3184
rect 3011 3144 3023 3184
rect 3031 3144 3043 3184
rect 3051 3144 3063 3172
rect 3071 3144 3083 3184
rect 3111 3144 3123 3184
rect 3131 3144 3143 3184
rect 3151 3144 3163 3172
rect 3171 3144 3183 3184
rect 3197 3144 3209 3184
rect 3217 3144 3229 3172
rect 3237 3144 3249 3184
rect 3257 3144 3269 3184
rect 3311 3144 3323 3184
rect 3331 3144 3343 3184
rect 3351 3144 3363 3172
rect 3371 3144 3383 3184
rect 3397 3144 3409 3184
rect 3417 3144 3429 3172
rect 3437 3144 3449 3184
rect 3457 3144 3469 3184
rect 3499 3144 3511 3184
rect 3529 3144 3541 3184
rect 3579 3144 3591 3184
rect 3609 3144 3621 3184
rect 3659 3144 3671 3184
rect 3689 3144 3701 3184
rect 3739 3144 3751 3184
rect 3769 3144 3781 3184
rect 3817 3144 3829 3164
rect 3839 3144 3851 3184
rect 3859 3144 3871 3184
rect 3919 3144 3931 3184
rect 3949 3144 3961 3184
rect 3991 3144 4003 3164
rect 4011 3144 4023 3164
rect 4031 3144 4043 3164
rect 4057 3144 4069 3164
rect 4079 3144 4091 3184
rect 4099 3144 4111 3184
rect 4151 3144 4163 3164
rect 4171 3144 4183 3164
rect 4211 3144 4223 3184
rect 4231 3144 4243 3184
rect 4251 3144 4263 3172
rect 4271 3144 4283 3184
rect 4311 3144 4323 3164
rect 4331 3144 4343 3164
rect 4357 3144 4369 3184
rect 4377 3144 4389 3172
rect 4397 3144 4409 3184
rect 4417 3144 4429 3184
rect 4479 3144 4491 3184
rect 4509 3144 4521 3184
rect 4541 3144 4553 3184
rect 4561 3144 4573 3164
rect 4593 3144 4605 3164
rect 4623 3144 4635 3164
rect 4645 3144 4657 3164
rect 4671 3144 4683 3164
rect 4699 3144 4711 3164
rect 4729 3144 4741 3164
rect 4751 3144 4763 3184
rect 52 3076 64 3116
rect 80 3076 92 3116
rect 108 3076 120 3116
rect 161 3076 173 3116
rect 181 3076 193 3116
rect 211 3076 223 3116
rect 237 3076 249 3116
rect 259 3096 271 3116
rect 289 3096 301 3116
rect 317 3096 329 3116
rect 343 3096 355 3116
rect 365 3096 377 3116
rect 395 3096 407 3116
rect 427 3096 439 3116
rect 447 3076 459 3116
rect 477 3076 489 3116
rect 497 3088 509 3116
rect 517 3076 529 3116
rect 537 3076 549 3116
rect 579 3076 591 3116
rect 609 3076 621 3116
rect 679 3076 691 3116
rect 709 3076 721 3116
rect 751 3096 763 3116
rect 771 3096 783 3116
rect 791 3096 803 3116
rect 819 3076 831 3116
rect 849 3076 861 3116
rect 911 3076 923 3116
rect 931 3076 943 3116
rect 951 3088 963 3116
rect 971 3076 983 3116
rect 1011 3076 1023 3116
rect 1031 3076 1043 3116
rect 1051 3088 1063 3116
rect 1071 3076 1083 3116
rect 1111 3096 1123 3116
rect 1131 3096 1143 3116
rect 1151 3096 1163 3116
rect 1191 3076 1203 3116
rect 1211 3076 1223 3116
rect 1231 3088 1243 3116
rect 1251 3076 1263 3116
rect 1279 3076 1291 3116
rect 1309 3076 1321 3116
rect 1371 3076 1383 3116
rect 1391 3076 1403 3116
rect 1419 3076 1431 3116
rect 1449 3076 1461 3116
rect 1499 3076 1511 3116
rect 1529 3076 1541 3116
rect 1577 3096 1589 3116
rect 1599 3076 1611 3116
rect 1619 3076 1631 3116
rect 1657 3076 1669 3116
rect 1677 3088 1689 3116
rect 1697 3076 1709 3116
rect 1717 3076 1729 3116
rect 1757 3076 1769 3116
rect 1777 3088 1789 3116
rect 1797 3076 1809 3116
rect 1817 3076 1829 3116
rect 1857 3096 1869 3116
rect 1877 3096 1889 3116
rect 1897 3096 1909 3116
rect 1940 3076 1952 3116
rect 1968 3076 1980 3116
rect 1990 3096 2002 3116
rect 2037 3096 2049 3116
rect 2057 3096 2069 3116
rect 2097 3076 2109 3116
rect 2117 3088 2129 3116
rect 2137 3076 2149 3116
rect 2157 3076 2169 3116
rect 2197 3096 2209 3116
rect 2217 3096 2229 3116
rect 2237 3096 2249 3116
rect 2299 3076 2311 3116
rect 2329 3076 2341 3116
rect 2357 3076 2369 3116
rect 2377 3088 2389 3116
rect 2397 3076 2409 3116
rect 2417 3076 2429 3116
rect 2457 3096 2469 3116
rect 2477 3096 2489 3116
rect 2517 3076 2529 3116
rect 2537 3088 2549 3116
rect 2557 3076 2569 3116
rect 2577 3076 2589 3116
rect 2617 3096 2629 3116
rect 2639 3076 2651 3116
rect 2659 3076 2671 3116
rect 2699 3076 2711 3116
rect 2729 3076 2741 3116
rect 2781 3076 2793 3116
rect 2801 3096 2813 3116
rect 2833 3096 2845 3116
rect 2863 3096 2875 3116
rect 2885 3096 2897 3116
rect 2911 3096 2923 3116
rect 2939 3096 2951 3116
rect 2969 3096 2981 3116
rect 2991 3076 3003 3116
rect 3031 3096 3043 3116
rect 3051 3096 3063 3116
rect 3071 3096 3083 3116
rect 3118 3096 3130 3116
rect 3140 3076 3152 3116
rect 3168 3076 3180 3116
rect 3197 3096 3209 3116
rect 3217 3096 3229 3116
rect 3237 3096 3249 3116
rect 3281 3076 3293 3116
rect 3301 3096 3313 3116
rect 3333 3096 3345 3116
rect 3363 3096 3375 3116
rect 3385 3096 3397 3116
rect 3411 3096 3423 3116
rect 3439 3096 3451 3116
rect 3469 3096 3481 3116
rect 3491 3076 3503 3116
rect 3521 3076 3533 3116
rect 3541 3096 3553 3116
rect 3573 3096 3585 3116
rect 3603 3096 3615 3116
rect 3625 3096 3637 3116
rect 3651 3096 3663 3116
rect 3679 3096 3691 3116
rect 3709 3096 3721 3116
rect 3731 3076 3743 3116
rect 3757 3096 3769 3116
rect 3777 3096 3789 3116
rect 3797 3096 3809 3116
rect 3851 3076 3863 3116
rect 3871 3076 3883 3116
rect 3891 3088 3903 3116
rect 3911 3076 3923 3116
rect 3951 3076 3963 3116
rect 3971 3076 3983 3116
rect 3991 3088 4003 3116
rect 4011 3076 4023 3116
rect 4037 3076 4049 3116
rect 4057 3088 4069 3116
rect 4077 3076 4089 3116
rect 4097 3076 4109 3116
rect 4137 3076 4149 3116
rect 4157 3088 4169 3116
rect 4177 3076 4189 3116
rect 4197 3076 4209 3116
rect 4237 3096 4249 3116
rect 4257 3096 4269 3116
rect 4298 3056 4310 3116
rect 4334 3058 4346 3116
rect 4397 3076 4409 3116
rect 4419 3096 4431 3116
rect 4449 3096 4461 3116
rect 4477 3096 4489 3116
rect 4503 3096 4515 3116
rect 4525 3096 4537 3116
rect 4555 3096 4567 3116
rect 4587 3096 4599 3116
rect 4607 3076 4619 3116
rect 4637 3076 4649 3116
rect 4657 3088 4669 3116
rect 4677 3076 4689 3116
rect 4697 3076 4709 3116
rect 31 2664 43 2684
rect 51 2664 63 2684
rect 91 2664 103 2704
rect 111 2664 123 2704
rect 131 2664 143 2692
rect 151 2664 163 2704
rect 180 2664 192 2704
rect 208 2664 220 2704
rect 236 2664 248 2704
rect 299 2664 311 2704
rect 329 2664 341 2704
rect 377 2664 389 2704
rect 407 2664 419 2704
rect 427 2664 439 2704
rect 491 2664 503 2704
rect 511 2664 523 2704
rect 531 2664 543 2692
rect 551 2664 563 2704
rect 579 2664 591 2704
rect 609 2664 621 2704
rect 671 2664 683 2704
rect 691 2664 703 2704
rect 731 2664 743 2704
rect 751 2664 763 2704
rect 779 2664 791 2704
rect 809 2664 821 2704
rect 857 2664 869 2704
rect 887 2664 899 2704
rect 907 2664 919 2704
rect 971 2664 983 2704
rect 991 2664 1003 2704
rect 1011 2664 1023 2692
rect 1031 2664 1043 2704
rect 1059 2664 1071 2704
rect 1089 2664 1101 2704
rect 1151 2664 1163 2704
rect 1171 2664 1183 2704
rect 1191 2664 1203 2692
rect 1211 2664 1223 2704
rect 1237 2664 1249 2704
rect 1259 2664 1271 2684
rect 1289 2664 1301 2684
rect 1317 2664 1329 2684
rect 1343 2664 1355 2684
rect 1365 2664 1377 2684
rect 1395 2664 1407 2684
rect 1427 2664 1439 2684
rect 1447 2664 1459 2704
rect 1489 2664 1501 2704
rect 1509 2664 1521 2704
rect 1531 2664 1543 2684
rect 1561 2664 1573 2704
rect 1581 2664 1593 2684
rect 1613 2664 1625 2684
rect 1643 2664 1655 2684
rect 1665 2664 1677 2684
rect 1691 2664 1703 2684
rect 1719 2664 1731 2684
rect 1749 2664 1761 2684
rect 1771 2664 1783 2704
rect 1797 2664 1809 2704
rect 1817 2664 1829 2692
rect 1837 2664 1849 2704
rect 1857 2664 1869 2704
rect 1897 2664 1909 2684
rect 1917 2664 1929 2684
rect 1957 2664 1969 2704
rect 1977 2664 1989 2694
rect 1997 2664 2009 2704
rect 2017 2676 2029 2704
rect 2037 2664 2049 2704
rect 2091 2664 2103 2684
rect 2111 2664 2123 2684
rect 2131 2664 2143 2684
rect 2171 2664 2183 2684
rect 2191 2664 2203 2684
rect 2211 2664 2223 2684
rect 2251 2664 2263 2684
rect 2271 2664 2283 2684
rect 2291 2664 2303 2684
rect 2317 2664 2329 2684
rect 2337 2664 2349 2684
rect 2391 2664 2403 2684
rect 2411 2664 2423 2684
rect 2431 2664 2443 2684
rect 2457 2664 2469 2684
rect 2477 2664 2489 2684
rect 2517 2664 2529 2704
rect 2547 2664 2559 2704
rect 2567 2664 2579 2704
rect 2617 2664 2629 2704
rect 2637 2664 2649 2692
rect 2657 2664 2669 2704
rect 2677 2664 2689 2704
rect 2717 2664 2729 2704
rect 2737 2664 2749 2692
rect 2757 2664 2769 2704
rect 2777 2664 2789 2704
rect 2819 2664 2831 2704
rect 2849 2664 2861 2704
rect 2901 2664 2913 2704
rect 2921 2664 2933 2684
rect 2953 2664 2965 2684
rect 2983 2664 2995 2684
rect 3005 2664 3017 2684
rect 3031 2664 3043 2684
rect 3059 2664 3071 2684
rect 3089 2664 3101 2684
rect 3111 2664 3123 2704
rect 3141 2664 3153 2704
rect 3161 2664 3173 2684
rect 3193 2664 3205 2684
rect 3223 2664 3235 2684
rect 3245 2664 3257 2684
rect 3271 2664 3283 2684
rect 3299 2664 3311 2684
rect 3329 2664 3341 2684
rect 3351 2664 3363 2704
rect 3391 2664 3403 2684
rect 3411 2664 3423 2684
rect 3451 2664 3463 2684
rect 3471 2664 3483 2684
rect 3491 2664 3503 2684
rect 3531 2664 3543 2704
rect 3551 2664 3563 2704
rect 3581 2664 3593 2704
rect 3601 2664 3613 2684
rect 3633 2664 3645 2684
rect 3663 2664 3675 2684
rect 3685 2664 3697 2684
rect 3711 2664 3723 2684
rect 3739 2664 3751 2684
rect 3769 2664 3781 2684
rect 3791 2664 3803 2704
rect 3852 2664 3864 2704
rect 3880 2664 3892 2704
rect 3908 2664 3920 2704
rect 3951 2664 3963 2684
rect 3971 2664 3983 2684
rect 3991 2664 4003 2684
rect 4017 2664 4029 2704
rect 4037 2664 4049 2692
rect 4057 2664 4069 2704
rect 4077 2664 4089 2704
rect 4131 2664 4143 2704
rect 4151 2664 4163 2704
rect 4171 2664 4183 2692
rect 4191 2664 4203 2704
rect 4217 2664 4229 2684
rect 4237 2664 4249 2684
rect 4257 2664 4269 2684
rect 4301 2664 4313 2704
rect 4321 2664 4333 2684
rect 4353 2664 4365 2684
rect 4383 2664 4395 2684
rect 4405 2664 4417 2684
rect 4431 2664 4443 2684
rect 4459 2664 4471 2684
rect 4489 2664 4501 2684
rect 4511 2664 4523 2704
rect 4537 2664 4549 2704
rect 4557 2664 4569 2692
rect 4577 2664 4589 2704
rect 4597 2664 4609 2704
rect 4639 2664 4651 2704
rect 4669 2664 4681 2704
rect 18 2576 30 2636
rect 54 2578 66 2636
rect 120 2596 132 2636
rect 148 2596 160 2636
rect 170 2616 182 2636
rect 231 2616 243 2636
rect 251 2616 263 2636
rect 301 2596 313 2636
rect 321 2596 333 2636
rect 351 2596 363 2636
rect 398 2616 410 2636
rect 420 2596 432 2636
rect 448 2596 460 2636
rect 514 2578 526 2636
rect 550 2576 562 2636
rect 591 2596 603 2636
rect 611 2596 623 2636
rect 631 2608 643 2636
rect 651 2596 663 2636
rect 691 2596 703 2636
rect 711 2596 723 2636
rect 759 2596 771 2636
rect 789 2596 801 2636
rect 854 2578 866 2636
rect 890 2576 902 2636
rect 931 2596 943 2636
rect 951 2596 963 2636
rect 971 2608 983 2636
rect 991 2596 1003 2636
rect 1019 2596 1031 2636
rect 1049 2596 1061 2636
rect 1134 2578 1146 2636
rect 1170 2576 1182 2636
rect 1211 2616 1223 2636
rect 1231 2616 1243 2636
rect 1271 2596 1283 2636
rect 1291 2596 1303 2636
rect 1311 2608 1323 2636
rect 1331 2596 1343 2636
rect 1359 2596 1371 2636
rect 1389 2596 1401 2636
rect 1437 2596 1449 2636
rect 1457 2596 1469 2636
rect 1519 2596 1531 2636
rect 1549 2596 1561 2636
rect 1581 2596 1593 2636
rect 1601 2616 1613 2636
rect 1633 2616 1645 2636
rect 1663 2616 1675 2636
rect 1685 2616 1697 2636
rect 1711 2616 1723 2636
rect 1739 2616 1751 2636
rect 1769 2616 1781 2636
rect 1791 2596 1803 2636
rect 1819 2596 1831 2636
rect 1849 2596 1861 2636
rect 1899 2596 1911 2636
rect 1929 2596 1941 2636
rect 1978 2576 1990 2636
rect 2014 2578 2026 2636
rect 2077 2616 2089 2636
rect 2097 2616 2109 2636
rect 2117 2616 2129 2636
rect 2171 2616 2183 2636
rect 2191 2616 2203 2636
rect 2231 2616 2243 2636
rect 2251 2616 2263 2636
rect 2271 2616 2283 2636
rect 2311 2616 2323 2636
rect 2331 2616 2343 2636
rect 2371 2596 2383 2636
rect 2391 2596 2403 2636
rect 2411 2608 2423 2636
rect 2431 2596 2443 2636
rect 2457 2616 2469 2636
rect 2477 2616 2489 2636
rect 2497 2616 2509 2636
rect 2537 2596 2549 2636
rect 2567 2596 2579 2636
rect 2587 2596 2599 2636
rect 2637 2596 2649 2636
rect 2657 2608 2669 2636
rect 2677 2596 2689 2636
rect 2697 2596 2709 2636
rect 2759 2596 2771 2636
rect 2789 2596 2801 2636
rect 2817 2616 2829 2636
rect 2837 2616 2849 2636
rect 2857 2616 2869 2636
rect 2877 2596 2889 2636
rect 2919 2596 2931 2636
rect 2949 2596 2961 2636
rect 2997 2616 3009 2636
rect 3019 2596 3031 2636
rect 3039 2596 3051 2636
rect 3077 2596 3089 2636
rect 3097 2608 3109 2636
rect 3117 2596 3129 2636
rect 3137 2596 3149 2636
rect 3189 2596 3201 2636
rect 3209 2596 3221 2636
rect 3231 2616 3243 2636
rect 3279 2596 3291 2636
rect 3309 2596 3321 2636
rect 3340 2596 3352 2636
rect 3368 2596 3380 2636
rect 3396 2596 3408 2636
rect 3457 2616 3469 2636
rect 3479 2596 3491 2636
rect 3499 2596 3511 2636
rect 3549 2596 3561 2636
rect 3569 2596 3581 2636
rect 3591 2616 3603 2636
rect 3621 2596 3633 2636
rect 3641 2616 3653 2636
rect 3673 2616 3685 2636
rect 3703 2616 3715 2636
rect 3725 2616 3737 2636
rect 3751 2616 3763 2636
rect 3779 2616 3791 2636
rect 3809 2616 3821 2636
rect 3831 2596 3843 2636
rect 3878 2616 3890 2636
rect 3900 2596 3912 2636
rect 3928 2596 3940 2636
rect 3957 2616 3969 2636
rect 3977 2616 3989 2636
rect 3997 2616 4009 2636
rect 4037 2596 4049 2636
rect 4057 2596 4069 2636
rect 4077 2596 4089 2636
rect 4097 2596 4109 2636
rect 4117 2596 4129 2636
rect 4137 2596 4149 2636
rect 4157 2596 4169 2636
rect 4177 2596 4189 2636
rect 4197 2596 4209 2636
rect 4241 2596 4253 2636
rect 4261 2616 4273 2636
rect 4293 2616 4305 2636
rect 4323 2616 4335 2636
rect 4345 2616 4357 2636
rect 4371 2616 4383 2636
rect 4399 2616 4411 2636
rect 4429 2616 4441 2636
rect 4451 2596 4463 2636
rect 4477 2596 4489 2636
rect 4497 2608 4509 2636
rect 4517 2596 4529 2636
rect 4537 2596 4549 2636
rect 4579 2596 4591 2636
rect 4609 2596 4621 2636
rect 4659 2596 4671 2636
rect 4689 2596 4701 2636
rect 54 2184 66 2242
rect 90 2184 102 2244
rect 131 2184 143 2224
rect 151 2184 163 2224
rect 171 2184 183 2212
rect 191 2184 203 2224
rect 217 2184 229 2224
rect 237 2184 249 2212
rect 257 2184 269 2224
rect 277 2184 289 2224
rect 318 2184 330 2244
rect 354 2184 366 2242
rect 420 2184 432 2224
rect 448 2184 460 2224
rect 470 2184 482 2204
rect 517 2184 529 2224
rect 537 2184 549 2212
rect 557 2184 569 2224
rect 577 2184 589 2224
rect 638 2184 650 2204
rect 660 2184 672 2224
rect 688 2184 700 2224
rect 717 2184 729 2204
rect 737 2184 749 2204
rect 801 2184 813 2224
rect 821 2184 833 2224
rect 851 2184 863 2224
rect 879 2184 891 2224
rect 909 2184 921 2224
rect 957 2184 969 2224
rect 987 2184 999 2224
rect 1007 2184 1019 2224
rect 1071 2184 1083 2224
rect 1091 2184 1103 2224
rect 1111 2184 1123 2212
rect 1131 2184 1143 2224
rect 1171 2184 1183 2224
rect 1191 2184 1203 2224
rect 1211 2184 1223 2212
rect 1231 2184 1243 2224
rect 1261 2184 1273 2224
rect 1281 2184 1293 2204
rect 1313 2184 1325 2204
rect 1343 2184 1355 2204
rect 1365 2184 1377 2204
rect 1391 2184 1403 2204
rect 1419 2184 1431 2204
rect 1449 2184 1461 2204
rect 1471 2184 1483 2224
rect 1511 2184 1523 2224
rect 1531 2184 1543 2224
rect 1551 2184 1563 2212
rect 1571 2184 1583 2224
rect 1601 2184 1613 2224
rect 1621 2184 1633 2204
rect 1653 2184 1665 2204
rect 1683 2184 1695 2204
rect 1705 2184 1717 2204
rect 1731 2184 1743 2204
rect 1759 2184 1771 2204
rect 1789 2184 1801 2204
rect 1811 2184 1823 2224
rect 1851 2184 1863 2204
rect 1871 2184 1883 2204
rect 1911 2184 1923 2204
rect 1931 2184 1943 2204
rect 1957 2184 1969 2224
rect 1977 2184 1989 2212
rect 1997 2184 2009 2224
rect 2017 2184 2029 2224
rect 2061 2184 2073 2224
rect 2081 2184 2093 2204
rect 2113 2184 2125 2204
rect 2143 2184 2155 2204
rect 2165 2184 2177 2204
rect 2191 2184 2203 2204
rect 2219 2184 2231 2204
rect 2249 2184 2261 2204
rect 2271 2184 2283 2224
rect 2318 2184 2330 2204
rect 2340 2184 2352 2224
rect 2368 2184 2380 2224
rect 2418 2184 2430 2204
rect 2440 2184 2452 2224
rect 2468 2184 2480 2224
rect 2498 2184 2510 2244
rect 2534 2184 2546 2242
rect 2597 2184 2609 2224
rect 2627 2184 2639 2224
rect 2647 2184 2659 2224
rect 2697 2184 2709 2224
rect 2719 2184 2731 2204
rect 2749 2184 2761 2204
rect 2777 2184 2789 2204
rect 2803 2184 2815 2204
rect 2825 2184 2837 2204
rect 2855 2184 2867 2204
rect 2887 2184 2899 2204
rect 2907 2184 2919 2224
rect 2951 2184 2963 2224
rect 2971 2184 2983 2224
rect 2991 2184 3003 2212
rect 3011 2184 3023 2224
rect 3051 2184 3063 2224
rect 3071 2184 3083 2224
rect 3091 2184 3103 2212
rect 3111 2184 3123 2224
rect 3137 2184 3149 2224
rect 3157 2184 3169 2212
rect 3177 2184 3189 2224
rect 3197 2184 3209 2224
rect 3237 2184 3249 2224
rect 3259 2184 3271 2204
rect 3289 2184 3301 2204
rect 3317 2184 3329 2204
rect 3343 2184 3355 2204
rect 3365 2184 3377 2204
rect 3395 2184 3407 2204
rect 3427 2184 3439 2204
rect 3447 2184 3459 2224
rect 3491 2184 3503 2224
rect 3511 2184 3523 2224
rect 3531 2184 3543 2212
rect 3551 2184 3563 2224
rect 3591 2184 3603 2204
rect 3611 2184 3623 2204
rect 3631 2184 3643 2204
rect 3657 2184 3669 2204
rect 3677 2184 3689 2204
rect 3697 2184 3709 2204
rect 3717 2184 3729 2224
rect 3779 2184 3791 2224
rect 3809 2184 3821 2224
rect 3872 2184 3884 2224
rect 3900 2184 3912 2224
rect 3928 2184 3940 2224
rect 3992 2184 4004 2224
rect 4020 2184 4032 2224
rect 4048 2184 4060 2224
rect 4081 2184 4093 2224
rect 4101 2184 4113 2204
rect 4133 2184 4145 2204
rect 4163 2184 4175 2204
rect 4185 2184 4197 2204
rect 4211 2184 4223 2204
rect 4239 2184 4251 2204
rect 4269 2184 4281 2204
rect 4291 2184 4303 2224
rect 4317 2184 4329 2224
rect 4339 2184 4351 2204
rect 4369 2184 4381 2204
rect 4397 2184 4409 2204
rect 4423 2184 4435 2204
rect 4445 2184 4457 2204
rect 4475 2184 4487 2204
rect 4507 2184 4519 2204
rect 4527 2184 4539 2224
rect 4557 2184 4569 2224
rect 4577 2184 4589 2212
rect 4597 2184 4609 2224
rect 4617 2184 4629 2224
rect 4659 2184 4671 2224
rect 4689 2184 4701 2224
rect 29 2116 41 2156
rect 49 2116 61 2156
rect 71 2136 83 2156
rect 111 2116 123 2156
rect 131 2116 143 2156
rect 151 2128 163 2156
rect 171 2116 183 2156
rect 234 2098 246 2156
rect 270 2096 282 2156
rect 300 2116 312 2156
rect 328 2116 340 2156
rect 350 2136 362 2156
rect 400 2116 412 2156
rect 428 2116 440 2156
rect 450 2136 462 2156
rect 498 2096 510 2156
rect 534 2098 546 2156
rect 598 2096 610 2156
rect 634 2098 646 2156
rect 700 2116 712 2156
rect 728 2116 740 2156
rect 750 2136 762 2156
rect 811 2116 823 2156
rect 831 2116 843 2156
rect 851 2128 863 2156
rect 871 2116 883 2156
rect 898 2096 910 2156
rect 934 2098 946 2156
rect 998 2096 1010 2156
rect 1034 2098 1046 2156
rect 1098 2096 1110 2156
rect 1134 2098 1146 2156
rect 1200 2116 1212 2156
rect 1228 2116 1240 2156
rect 1250 2136 1262 2156
rect 1297 2136 1309 2156
rect 1317 2136 1329 2156
rect 1337 2136 1349 2156
rect 1399 2116 1411 2156
rect 1429 2116 1441 2156
rect 1479 2116 1491 2156
rect 1509 2116 1521 2156
rect 1539 2116 1551 2156
rect 1569 2116 1581 2156
rect 1631 2116 1643 2156
rect 1651 2116 1663 2156
rect 1671 2128 1683 2156
rect 1691 2116 1703 2156
rect 1720 2116 1732 2156
rect 1748 2116 1760 2156
rect 1770 2136 1782 2156
rect 1817 2136 1829 2156
rect 1837 2136 1849 2156
rect 1857 2136 1869 2156
rect 1911 2116 1923 2156
rect 1931 2116 1943 2156
rect 1951 2128 1963 2156
rect 1971 2116 1983 2156
rect 1997 2116 2009 2156
rect 2017 2128 2029 2156
rect 2037 2116 2049 2156
rect 2057 2116 2069 2156
rect 2111 2116 2123 2156
rect 2131 2116 2143 2156
rect 2151 2128 2163 2156
rect 2171 2116 2183 2156
rect 2211 2116 2223 2156
rect 2231 2116 2243 2156
rect 2251 2116 2263 2156
rect 2271 2116 2283 2156
rect 2291 2116 2303 2156
rect 2311 2116 2323 2156
rect 2331 2116 2343 2156
rect 2351 2116 2363 2156
rect 2371 2116 2383 2156
rect 2399 2116 2411 2156
rect 2429 2116 2441 2156
rect 2501 2116 2513 2156
rect 2521 2116 2533 2156
rect 2551 2116 2563 2156
rect 2577 2136 2589 2156
rect 2597 2136 2609 2156
rect 2617 2136 2629 2156
rect 2637 2116 2649 2156
rect 2699 2116 2711 2156
rect 2729 2116 2741 2156
rect 2759 2116 2771 2156
rect 2789 2116 2801 2156
rect 2841 2116 2853 2156
rect 2861 2136 2873 2156
rect 2893 2136 2905 2156
rect 2923 2136 2935 2156
rect 2945 2136 2957 2156
rect 2971 2136 2983 2156
rect 2999 2136 3011 2156
rect 3029 2136 3041 2156
rect 3051 2116 3063 2156
rect 3098 2136 3110 2156
rect 3120 2116 3132 2156
rect 3148 2116 3160 2156
rect 3177 2136 3189 2156
rect 3197 2136 3209 2156
rect 3217 2136 3229 2156
rect 3292 2116 3304 2156
rect 3320 2116 3332 2156
rect 3348 2116 3360 2156
rect 3381 2116 3393 2156
rect 3401 2136 3413 2156
rect 3433 2136 3445 2156
rect 3463 2136 3475 2156
rect 3485 2136 3497 2156
rect 3511 2136 3523 2156
rect 3539 2136 3551 2156
rect 3569 2136 3581 2156
rect 3591 2116 3603 2156
rect 3617 2116 3629 2156
rect 3637 2128 3649 2156
rect 3657 2116 3669 2156
rect 3677 2116 3689 2156
rect 3721 2116 3733 2156
rect 3741 2136 3753 2156
rect 3773 2136 3785 2156
rect 3803 2136 3815 2156
rect 3825 2136 3837 2156
rect 3851 2136 3863 2156
rect 3879 2136 3891 2156
rect 3909 2136 3921 2156
rect 3931 2116 3943 2156
rect 3957 2116 3969 2156
rect 3979 2136 3991 2156
rect 4009 2136 4021 2156
rect 4037 2136 4049 2156
rect 4063 2136 4075 2156
rect 4085 2136 4097 2156
rect 4115 2136 4127 2156
rect 4147 2136 4159 2156
rect 4167 2116 4179 2156
rect 4232 2116 4244 2156
rect 4260 2116 4272 2156
rect 4288 2116 4300 2156
rect 4317 2136 4329 2156
rect 4337 2136 4349 2156
rect 4391 2136 4403 2156
rect 4411 2136 4423 2156
rect 4431 2136 4443 2156
rect 4471 2136 4483 2156
rect 4491 2136 4503 2156
rect 4511 2136 4523 2156
rect 4537 2116 4549 2156
rect 4559 2136 4571 2156
rect 4589 2136 4601 2156
rect 4617 2136 4629 2156
rect 4643 2136 4655 2156
rect 4665 2136 4677 2156
rect 4695 2136 4707 2156
rect 4727 2136 4739 2156
rect 4747 2116 4759 2156
rect 52 1704 64 1744
rect 80 1704 92 1744
rect 108 1704 120 1744
rect 137 1704 149 1744
rect 157 1704 169 1732
rect 177 1704 189 1744
rect 197 1704 209 1744
rect 239 1704 251 1744
rect 269 1704 281 1744
rect 354 1704 366 1762
rect 390 1704 402 1764
rect 420 1704 432 1744
rect 448 1704 460 1744
rect 476 1704 488 1744
rect 537 1704 549 1744
rect 567 1704 579 1744
rect 587 1704 599 1744
rect 651 1704 663 1744
rect 671 1704 683 1744
rect 697 1704 709 1724
rect 719 1704 731 1744
rect 739 1704 751 1744
rect 791 1704 803 1744
rect 811 1704 823 1744
rect 831 1704 843 1732
rect 851 1704 863 1744
rect 877 1704 889 1744
rect 897 1704 909 1732
rect 917 1704 929 1744
rect 937 1704 949 1744
rect 978 1704 990 1764
rect 1014 1704 1026 1762
rect 1077 1704 1089 1724
rect 1097 1704 1109 1724
rect 1138 1704 1150 1764
rect 1174 1704 1186 1762
rect 1238 1704 1250 1764
rect 1274 1704 1286 1762
rect 1351 1704 1363 1724
rect 1371 1704 1383 1724
rect 1432 1704 1444 1744
rect 1460 1704 1472 1744
rect 1488 1704 1500 1744
rect 1518 1704 1530 1764
rect 1554 1704 1566 1762
rect 1617 1704 1629 1724
rect 1637 1704 1649 1724
rect 1691 1704 1703 1744
rect 1711 1704 1723 1744
rect 1774 1704 1786 1762
rect 1810 1704 1822 1764
rect 1837 1704 1849 1744
rect 1867 1704 1879 1744
rect 1887 1704 1899 1744
rect 1941 1704 1953 1744
rect 1961 1704 1973 1724
rect 1993 1704 2005 1724
rect 2023 1704 2035 1724
rect 2045 1704 2057 1724
rect 2071 1704 2083 1724
rect 2099 1704 2111 1724
rect 2129 1704 2141 1724
rect 2151 1704 2163 1744
rect 2191 1704 2203 1724
rect 2211 1704 2223 1724
rect 2231 1704 2243 1724
rect 2257 1704 2269 1724
rect 2277 1704 2289 1724
rect 2317 1704 2329 1744
rect 2337 1704 2349 1732
rect 2357 1704 2369 1744
rect 2377 1704 2389 1744
rect 2417 1704 2429 1724
rect 2437 1704 2449 1724
rect 2457 1704 2469 1724
rect 2497 1704 2509 1724
rect 2517 1704 2529 1724
rect 2537 1704 2549 1724
rect 2577 1704 2589 1744
rect 2597 1704 2609 1732
rect 2617 1704 2629 1744
rect 2637 1704 2649 1744
rect 2699 1704 2711 1744
rect 2729 1704 2741 1744
rect 2771 1704 2783 1724
rect 2791 1704 2803 1724
rect 2811 1704 2823 1724
rect 2837 1704 2849 1744
rect 2857 1704 2869 1732
rect 2877 1704 2889 1744
rect 2897 1704 2909 1744
rect 2937 1704 2949 1724
rect 2957 1704 2969 1724
rect 3011 1704 3023 1724
rect 3031 1704 3043 1724
rect 3051 1704 3063 1724
rect 3077 1704 3089 1744
rect 3099 1704 3111 1724
rect 3129 1704 3141 1724
rect 3157 1704 3169 1724
rect 3183 1704 3195 1724
rect 3205 1704 3217 1724
rect 3235 1704 3247 1724
rect 3267 1704 3279 1724
rect 3287 1704 3299 1744
rect 3317 1704 3329 1744
rect 3337 1704 3349 1732
rect 3357 1704 3369 1744
rect 3377 1704 3389 1744
rect 3419 1704 3431 1744
rect 3449 1704 3461 1744
rect 3497 1704 3509 1744
rect 3519 1704 3531 1724
rect 3549 1704 3561 1724
rect 3577 1704 3589 1724
rect 3603 1704 3615 1724
rect 3625 1704 3637 1724
rect 3655 1704 3667 1724
rect 3687 1704 3699 1724
rect 3707 1704 3719 1744
rect 3737 1704 3749 1724
rect 3759 1704 3771 1744
rect 3779 1704 3791 1744
rect 3839 1704 3851 1744
rect 3869 1704 3881 1744
rect 3911 1704 3923 1744
rect 3931 1704 3943 1744
rect 3951 1704 3963 1732
rect 3971 1704 3983 1744
rect 4011 1704 4023 1744
rect 4031 1704 4043 1744
rect 4051 1704 4063 1732
rect 4071 1704 4083 1744
rect 4097 1704 4109 1724
rect 4117 1704 4129 1724
rect 4137 1704 4149 1724
rect 4157 1704 4169 1744
rect 4211 1704 4223 1724
rect 4231 1704 4243 1724
rect 4260 1704 4272 1744
rect 4288 1704 4300 1744
rect 4310 1704 4322 1724
rect 4371 1704 4383 1724
rect 4391 1704 4403 1724
rect 4411 1704 4423 1724
rect 4437 1704 4449 1744
rect 4459 1704 4471 1724
rect 4489 1704 4501 1724
rect 4517 1704 4529 1724
rect 4543 1704 4555 1724
rect 4565 1704 4577 1724
rect 4595 1704 4607 1724
rect 4627 1704 4639 1724
rect 4647 1704 4659 1744
rect 4699 1704 4711 1744
rect 4729 1704 4741 1744
rect 31 1656 43 1676
rect 51 1656 63 1676
rect 98 1656 110 1676
rect 120 1636 132 1676
rect 148 1636 160 1676
rect 178 1616 190 1676
rect 214 1618 226 1676
rect 279 1636 291 1676
rect 309 1636 321 1676
rect 371 1636 383 1676
rect 391 1636 403 1676
rect 411 1648 423 1676
rect 431 1636 443 1676
rect 469 1636 481 1676
rect 489 1636 501 1676
rect 511 1656 523 1676
rect 551 1656 563 1676
rect 571 1656 583 1676
rect 598 1616 610 1676
rect 634 1618 646 1676
rect 700 1636 712 1676
rect 728 1636 740 1676
rect 750 1656 762 1676
rect 798 1616 810 1676
rect 834 1618 846 1676
rect 900 1636 912 1676
rect 928 1636 940 1676
rect 950 1656 962 1676
rect 998 1616 1010 1676
rect 1034 1618 1046 1676
rect 1111 1636 1123 1676
rect 1131 1636 1143 1676
rect 1151 1648 1163 1676
rect 1171 1636 1183 1676
rect 1198 1616 1210 1676
rect 1234 1618 1246 1676
rect 1300 1636 1312 1676
rect 1328 1636 1340 1676
rect 1350 1656 1362 1676
rect 1411 1656 1423 1676
rect 1431 1656 1443 1676
rect 1458 1616 1470 1676
rect 1494 1618 1506 1676
rect 1560 1636 1572 1676
rect 1588 1636 1600 1676
rect 1610 1656 1622 1676
rect 1658 1616 1670 1676
rect 1694 1618 1706 1676
rect 1757 1636 1769 1676
rect 1777 1648 1789 1676
rect 1797 1636 1809 1676
rect 1817 1636 1829 1676
rect 1878 1656 1890 1676
rect 1900 1636 1912 1676
rect 1928 1636 1940 1676
rect 1957 1656 1969 1676
rect 1977 1656 1989 1676
rect 2018 1616 2030 1676
rect 2054 1618 2066 1676
rect 2131 1636 2143 1676
rect 2151 1636 2163 1676
rect 2171 1648 2183 1676
rect 2191 1636 2203 1676
rect 2217 1656 2229 1676
rect 2237 1656 2249 1676
rect 2277 1636 2289 1676
rect 2299 1656 2311 1676
rect 2329 1656 2341 1676
rect 2357 1656 2369 1676
rect 2383 1656 2395 1676
rect 2405 1656 2417 1676
rect 2435 1656 2447 1676
rect 2467 1656 2479 1676
rect 2487 1636 2499 1676
rect 2531 1636 2543 1676
rect 2551 1636 2563 1676
rect 2571 1648 2583 1676
rect 2591 1636 2603 1676
rect 2641 1636 2653 1676
rect 2661 1636 2673 1676
rect 2691 1636 2703 1676
rect 2717 1656 2729 1676
rect 2737 1656 2749 1676
rect 2757 1656 2769 1676
rect 2800 1636 2812 1676
rect 2828 1636 2840 1676
rect 2850 1656 2862 1676
rect 2911 1656 2923 1676
rect 2931 1656 2943 1676
rect 2951 1656 2963 1676
rect 2991 1656 3003 1676
rect 3011 1656 3023 1676
rect 3051 1656 3063 1676
rect 3071 1656 3083 1676
rect 3097 1636 3109 1676
rect 3117 1648 3129 1676
rect 3137 1636 3149 1676
rect 3157 1636 3169 1676
rect 3199 1636 3211 1676
rect 3229 1636 3241 1676
rect 3299 1636 3311 1676
rect 3329 1636 3341 1676
rect 3371 1636 3383 1676
rect 3391 1636 3403 1676
rect 3411 1648 3423 1676
rect 3431 1636 3443 1676
rect 3461 1636 3473 1676
rect 3481 1656 3493 1676
rect 3513 1656 3525 1676
rect 3543 1656 3555 1676
rect 3565 1656 3577 1676
rect 3591 1656 3603 1676
rect 3619 1656 3631 1676
rect 3649 1656 3661 1676
rect 3671 1636 3683 1676
rect 3697 1656 3709 1676
rect 3717 1656 3729 1676
rect 3771 1656 3783 1676
rect 3791 1656 3803 1676
rect 3831 1636 3843 1676
rect 3851 1636 3863 1676
rect 3871 1648 3883 1676
rect 3891 1636 3903 1676
rect 3917 1656 3929 1676
rect 3937 1656 3949 1676
rect 3957 1656 3969 1676
rect 3997 1656 4009 1676
rect 4017 1656 4029 1676
rect 4037 1656 4049 1676
rect 4077 1656 4089 1676
rect 4097 1656 4109 1676
rect 4140 1636 4152 1676
rect 4168 1636 4180 1676
rect 4190 1656 4202 1676
rect 4237 1656 4249 1676
rect 4257 1656 4269 1676
rect 4277 1656 4289 1676
rect 4320 1636 4332 1676
rect 4348 1636 4360 1676
rect 4370 1656 4382 1676
rect 4417 1656 4429 1676
rect 4437 1656 4449 1676
rect 4477 1656 4489 1676
rect 4497 1656 4509 1676
rect 4551 1656 4563 1676
rect 4571 1656 4583 1676
rect 4597 1636 4609 1676
rect 4617 1648 4629 1676
rect 4637 1636 4649 1676
rect 4657 1636 4669 1676
rect 4699 1636 4711 1676
rect 4729 1636 4741 1676
rect 38 1224 50 1244
rect 60 1224 72 1264
rect 88 1224 100 1264
rect 118 1224 130 1284
rect 154 1224 166 1282
rect 218 1224 230 1284
rect 254 1224 266 1282
rect 339 1224 351 1264
rect 369 1224 381 1264
rect 397 1224 409 1264
rect 417 1224 429 1252
rect 437 1224 449 1264
rect 457 1224 469 1264
rect 500 1224 512 1264
rect 528 1224 540 1264
rect 550 1224 562 1244
rect 597 1224 609 1264
rect 617 1224 629 1252
rect 637 1224 649 1264
rect 657 1224 669 1264
rect 697 1224 709 1264
rect 717 1224 729 1252
rect 737 1224 749 1264
rect 757 1224 769 1264
rect 797 1224 809 1264
rect 827 1224 839 1264
rect 847 1224 859 1264
rect 919 1224 931 1264
rect 949 1224 961 1264
rect 979 1224 991 1264
rect 1009 1224 1021 1264
rect 1094 1224 1106 1282
rect 1130 1224 1142 1284
rect 1171 1224 1183 1244
rect 1191 1224 1203 1244
rect 1241 1224 1253 1264
rect 1261 1224 1273 1264
rect 1291 1224 1303 1264
rect 1317 1224 1329 1264
rect 1337 1224 1349 1252
rect 1357 1224 1369 1264
rect 1377 1224 1389 1264
rect 1431 1224 1443 1264
rect 1451 1224 1463 1264
rect 1471 1224 1483 1252
rect 1491 1224 1503 1264
rect 1519 1224 1531 1264
rect 1549 1224 1561 1264
rect 1597 1224 1609 1264
rect 1617 1224 1629 1252
rect 1637 1224 1649 1264
rect 1657 1224 1669 1264
rect 1699 1224 1711 1264
rect 1729 1224 1741 1264
rect 1780 1224 1792 1264
rect 1808 1224 1820 1264
rect 1830 1224 1842 1244
rect 1878 1224 1890 1284
rect 1914 1224 1926 1282
rect 1977 1224 1989 1264
rect 1997 1224 2009 1252
rect 2017 1224 2029 1264
rect 2037 1224 2049 1264
rect 2077 1224 2089 1244
rect 2097 1224 2109 1244
rect 2138 1224 2150 1284
rect 2174 1224 2186 1282
rect 2239 1224 2251 1264
rect 2269 1224 2281 1264
rect 2317 1224 2329 1244
rect 2337 1224 2349 1244
rect 2357 1224 2369 1244
rect 2377 1224 2389 1264
rect 2439 1224 2451 1264
rect 2469 1224 2481 1264
rect 2497 1224 2509 1244
rect 2517 1224 2529 1244
rect 2569 1224 2581 1264
rect 2589 1224 2601 1264
rect 2611 1224 2623 1244
rect 2637 1224 2649 1264
rect 2657 1224 2669 1252
rect 2677 1224 2689 1264
rect 2697 1224 2709 1264
rect 2751 1224 2763 1264
rect 2771 1236 2783 1264
rect 2791 1224 2803 1264
rect 2811 1224 2823 1254
rect 2831 1224 2843 1264
rect 2861 1224 2873 1264
rect 2881 1224 2893 1244
rect 2913 1224 2925 1244
rect 2943 1224 2955 1244
rect 2965 1224 2977 1244
rect 2991 1224 3003 1244
rect 3019 1224 3031 1244
rect 3049 1224 3061 1244
rect 3071 1224 3083 1264
rect 3111 1224 3123 1244
rect 3131 1224 3143 1244
rect 3151 1224 3163 1244
rect 3198 1224 3210 1244
rect 3220 1224 3232 1264
rect 3248 1224 3260 1264
rect 3281 1224 3293 1264
rect 3301 1224 3313 1244
rect 3333 1224 3345 1244
rect 3363 1224 3375 1244
rect 3385 1224 3397 1244
rect 3411 1224 3423 1244
rect 3439 1224 3451 1244
rect 3469 1224 3481 1244
rect 3491 1224 3503 1264
rect 3531 1224 3543 1244
rect 3551 1224 3563 1244
rect 3591 1224 3603 1244
rect 3611 1224 3623 1244
rect 3631 1224 3643 1244
rect 3671 1224 3683 1244
rect 3691 1224 3703 1244
rect 3711 1224 3723 1244
rect 3737 1224 3749 1244
rect 3757 1224 3769 1244
rect 3797 1224 3809 1264
rect 3819 1224 3831 1244
rect 3849 1224 3861 1244
rect 3877 1224 3889 1244
rect 3903 1224 3915 1244
rect 3925 1224 3937 1244
rect 3955 1224 3967 1244
rect 3987 1224 3999 1244
rect 4007 1224 4019 1264
rect 4037 1224 4049 1264
rect 4057 1224 4069 1252
rect 4077 1224 4089 1264
rect 4097 1224 4109 1264
rect 4139 1224 4151 1264
rect 4169 1224 4181 1264
rect 4229 1224 4241 1264
rect 4249 1224 4261 1264
rect 4271 1224 4283 1244
rect 4319 1224 4331 1264
rect 4349 1224 4361 1264
rect 4391 1224 4403 1264
rect 4411 1224 4423 1264
rect 4431 1224 4443 1252
rect 4451 1224 4463 1264
rect 4491 1224 4503 1264
rect 4511 1224 4523 1264
rect 4531 1224 4543 1252
rect 4551 1224 4563 1264
rect 4577 1224 4589 1244
rect 4597 1224 4609 1244
rect 4617 1224 4629 1244
rect 4657 1224 4669 1244
rect 4677 1224 4689 1244
rect 4731 1224 4743 1244
rect 4751 1224 4763 1244
rect 31 1156 43 1196
rect 51 1156 63 1196
rect 71 1168 83 1196
rect 91 1156 103 1196
rect 117 1156 129 1196
rect 137 1168 149 1196
rect 157 1156 169 1196
rect 177 1156 189 1196
rect 218 1136 230 1196
rect 254 1138 266 1196
rect 320 1156 332 1196
rect 348 1156 360 1196
rect 370 1176 382 1196
rect 418 1136 430 1196
rect 454 1138 466 1196
rect 520 1156 532 1196
rect 548 1156 560 1196
rect 570 1176 582 1196
rect 639 1156 651 1196
rect 669 1156 681 1196
rect 721 1156 733 1196
rect 741 1156 753 1196
rect 771 1156 783 1196
rect 834 1138 846 1196
rect 870 1136 882 1196
rect 911 1156 923 1196
rect 931 1156 943 1196
rect 951 1168 963 1196
rect 971 1156 983 1196
rect 997 1156 1009 1196
rect 1017 1168 1029 1196
rect 1037 1156 1049 1196
rect 1057 1156 1069 1196
rect 1111 1156 1123 1196
rect 1131 1156 1143 1196
rect 1151 1168 1163 1196
rect 1171 1156 1183 1196
rect 1219 1156 1231 1196
rect 1249 1156 1261 1196
rect 1301 1156 1313 1196
rect 1321 1156 1333 1196
rect 1351 1156 1363 1196
rect 1379 1156 1391 1196
rect 1409 1156 1421 1196
rect 1471 1156 1483 1196
rect 1491 1156 1503 1196
rect 1539 1156 1551 1196
rect 1569 1156 1581 1196
rect 1619 1156 1631 1196
rect 1649 1156 1661 1196
rect 1678 1136 1690 1196
rect 1714 1138 1726 1196
rect 1799 1156 1811 1196
rect 1829 1156 1841 1196
rect 1858 1136 1870 1196
rect 1894 1138 1906 1196
rect 1959 1156 1971 1196
rect 1989 1156 2001 1196
rect 2072 1156 2084 1196
rect 2100 1156 2112 1196
rect 2128 1156 2140 1196
rect 2194 1138 2206 1196
rect 2230 1136 2242 1196
rect 2279 1156 2291 1196
rect 2309 1156 2321 1196
rect 2340 1156 2352 1196
rect 2368 1156 2380 1196
rect 2390 1176 2402 1196
rect 2451 1176 2463 1196
rect 2471 1176 2483 1196
rect 2519 1156 2531 1196
rect 2549 1156 2561 1196
rect 2591 1156 2603 1196
rect 2611 1156 2623 1184
rect 2631 1156 2643 1196
rect 2651 1166 2663 1196
rect 2671 1156 2683 1196
rect 2697 1176 2709 1196
rect 2719 1156 2731 1196
rect 2739 1156 2751 1196
rect 2781 1156 2793 1196
rect 2801 1176 2813 1196
rect 2833 1176 2845 1196
rect 2863 1176 2875 1196
rect 2885 1176 2897 1196
rect 2911 1176 2923 1196
rect 2939 1176 2951 1196
rect 2969 1176 2981 1196
rect 2991 1156 3003 1196
rect 3019 1156 3031 1196
rect 3049 1156 3061 1196
rect 3111 1156 3123 1196
rect 3131 1156 3143 1196
rect 3151 1168 3163 1196
rect 3171 1156 3183 1196
rect 3197 1156 3209 1196
rect 3217 1156 3229 1196
rect 3237 1156 3249 1196
rect 3257 1156 3269 1196
rect 3277 1156 3289 1196
rect 3329 1156 3341 1196
rect 3349 1156 3361 1196
rect 3371 1176 3383 1196
rect 3397 1176 3409 1196
rect 3419 1156 3431 1196
rect 3439 1156 3451 1196
rect 3477 1156 3489 1196
rect 3497 1156 3509 1196
rect 3517 1156 3529 1196
rect 3537 1156 3549 1196
rect 3557 1156 3569 1196
rect 3577 1156 3589 1196
rect 3597 1156 3609 1196
rect 3617 1156 3629 1196
rect 3637 1156 3649 1196
rect 3677 1156 3689 1196
rect 3697 1156 3709 1196
rect 3717 1156 3729 1196
rect 3737 1156 3749 1196
rect 3757 1156 3769 1196
rect 3777 1156 3789 1196
rect 3797 1156 3809 1196
rect 3817 1156 3829 1196
rect 3837 1156 3849 1196
rect 3877 1176 3889 1196
rect 3899 1156 3911 1196
rect 3919 1156 3931 1196
rect 3959 1156 3971 1196
rect 3989 1156 4001 1196
rect 4037 1156 4049 1196
rect 4059 1176 4071 1196
rect 4089 1176 4101 1196
rect 4117 1176 4129 1196
rect 4143 1176 4155 1196
rect 4165 1176 4177 1196
rect 4195 1176 4207 1196
rect 4227 1176 4239 1196
rect 4247 1156 4259 1196
rect 4279 1156 4291 1196
rect 4309 1156 4321 1196
rect 4357 1156 4369 1196
rect 4377 1168 4389 1196
rect 4397 1156 4409 1196
rect 4417 1156 4429 1196
rect 4479 1156 4491 1196
rect 4509 1156 4521 1196
rect 4537 1156 4549 1196
rect 4557 1168 4569 1196
rect 4577 1156 4589 1196
rect 4597 1156 4609 1196
rect 4638 1136 4650 1196
rect 4674 1138 4686 1196
rect 39 744 51 784
rect 69 744 81 784
rect 121 744 133 784
rect 141 744 153 784
rect 171 744 183 784
rect 211 744 223 784
rect 231 744 243 784
rect 251 744 263 772
rect 271 744 283 784
rect 332 744 344 784
rect 360 744 372 784
rect 388 744 400 784
rect 429 744 441 784
rect 449 744 461 784
rect 471 744 483 764
rect 497 744 509 764
rect 517 744 529 764
rect 571 744 583 764
rect 591 744 603 764
rect 638 744 650 764
rect 660 744 672 784
rect 688 744 700 784
rect 718 744 730 804
rect 754 744 766 802
rect 841 744 853 784
rect 861 744 873 784
rect 891 744 903 784
rect 919 744 931 784
rect 949 744 961 784
rect 1034 744 1046 802
rect 1070 744 1082 804
rect 1097 744 1109 784
rect 1117 744 1129 772
rect 1137 744 1149 784
rect 1157 744 1169 784
rect 1234 744 1246 802
rect 1270 744 1282 804
rect 1297 744 1309 764
rect 1317 744 1329 764
rect 1357 744 1369 784
rect 1377 744 1389 772
rect 1397 744 1409 784
rect 1417 744 1429 784
rect 1479 744 1491 784
rect 1509 744 1521 784
rect 1539 744 1551 784
rect 1569 744 1581 784
rect 1631 744 1643 784
rect 1651 744 1663 784
rect 1671 744 1683 772
rect 1691 744 1703 784
rect 1717 744 1729 784
rect 1747 744 1759 784
rect 1767 744 1779 784
rect 1831 744 1843 764
rect 1851 744 1863 764
rect 1899 744 1911 784
rect 1929 744 1941 784
rect 1957 744 1969 764
rect 1977 744 1989 764
rect 2054 744 2066 802
rect 2090 744 2102 804
rect 2117 744 2129 764
rect 2137 744 2149 764
rect 2177 744 2189 784
rect 2197 744 2209 772
rect 2217 744 2229 784
rect 2237 744 2249 784
rect 2298 744 2310 764
rect 2320 744 2332 784
rect 2348 744 2360 784
rect 2377 744 2389 764
rect 2397 744 2409 764
rect 2438 744 2450 804
rect 2474 744 2486 802
rect 2574 744 2586 802
rect 2610 744 2622 804
rect 2640 744 2652 784
rect 2668 744 2680 784
rect 2690 744 2702 764
rect 2759 744 2771 784
rect 2789 744 2801 784
rect 2831 744 2843 784
rect 2851 756 2863 784
rect 2871 744 2883 784
rect 2891 744 2903 774
rect 2911 744 2923 784
rect 2951 744 2963 764
rect 2971 744 2983 764
rect 3011 744 3023 764
rect 3031 744 3043 764
rect 3051 744 3063 764
rect 3091 744 3103 764
rect 3111 744 3123 764
rect 3131 744 3143 764
rect 3157 744 3169 764
rect 3177 744 3189 764
rect 3217 744 3229 784
rect 3237 744 3249 772
rect 3257 744 3269 784
rect 3277 744 3289 784
rect 3319 744 3331 784
rect 3349 744 3361 784
rect 3397 744 3409 784
rect 3419 744 3431 764
rect 3449 744 3461 764
rect 3477 744 3489 764
rect 3503 744 3515 764
rect 3525 744 3537 764
rect 3555 744 3567 764
rect 3587 744 3599 764
rect 3607 744 3619 784
rect 3637 744 3649 764
rect 3659 744 3671 784
rect 3679 744 3691 784
rect 3721 744 3733 784
rect 3741 744 3753 764
rect 3773 744 3785 764
rect 3803 744 3815 764
rect 3825 744 3837 764
rect 3851 744 3863 764
rect 3879 744 3891 764
rect 3909 744 3921 764
rect 3931 744 3943 784
rect 3971 744 3983 784
rect 3991 744 4003 784
rect 4011 744 4023 772
rect 4031 744 4043 784
rect 4057 744 4069 784
rect 4079 744 4091 764
rect 4109 744 4121 764
rect 4137 744 4149 764
rect 4163 744 4175 764
rect 4185 744 4197 764
rect 4215 744 4227 764
rect 4247 744 4259 764
rect 4267 744 4279 784
rect 4301 744 4313 784
rect 4321 744 4333 764
rect 4353 744 4365 764
rect 4383 744 4395 764
rect 4405 744 4417 764
rect 4431 744 4443 764
rect 4459 744 4471 764
rect 4489 744 4501 764
rect 4511 744 4523 784
rect 4537 744 4549 784
rect 4557 744 4569 772
rect 4577 744 4589 784
rect 4597 744 4609 784
rect 4637 744 4649 784
rect 4657 744 4669 772
rect 4677 744 4689 784
rect 4697 744 4709 784
rect 31 696 43 716
rect 51 696 63 716
rect 71 696 83 716
rect 118 696 130 716
rect 140 676 152 716
rect 168 676 180 716
rect 197 696 209 716
rect 217 696 229 716
rect 278 696 290 716
rect 300 676 312 716
rect 328 676 340 716
rect 358 656 370 716
rect 394 658 406 716
rect 471 676 483 716
rect 491 676 503 716
rect 511 688 523 716
rect 531 676 543 716
rect 569 676 581 716
rect 589 676 601 716
rect 611 696 623 716
rect 651 676 663 716
rect 671 676 683 716
rect 691 688 703 716
rect 711 676 723 716
rect 749 676 761 716
rect 769 676 781 716
rect 791 696 803 716
rect 817 676 829 716
rect 847 676 859 716
rect 867 676 879 716
rect 917 676 929 716
rect 937 688 949 716
rect 957 676 969 716
rect 977 676 989 716
rect 1031 676 1043 716
rect 1051 676 1063 716
rect 1071 688 1083 716
rect 1091 676 1103 716
rect 1131 676 1143 716
rect 1151 676 1163 716
rect 1180 676 1192 716
rect 1208 676 1220 716
rect 1230 696 1242 716
rect 1291 696 1303 716
rect 1311 696 1323 716
rect 1337 676 1349 716
rect 1357 688 1369 716
rect 1377 676 1389 716
rect 1397 676 1409 716
rect 1437 676 1449 716
rect 1457 688 1469 716
rect 1477 676 1489 716
rect 1497 676 1509 716
rect 1558 696 1570 716
rect 1580 676 1592 716
rect 1608 676 1620 716
rect 1640 676 1652 716
rect 1668 676 1680 716
rect 1690 696 1702 716
rect 1738 656 1750 716
rect 1774 658 1786 716
rect 1837 676 1849 716
rect 1857 688 1869 716
rect 1877 676 1889 716
rect 1897 676 1909 716
rect 1958 696 1970 716
rect 1980 676 1992 716
rect 2008 676 2020 716
rect 2037 676 2049 716
rect 2057 688 2069 716
rect 2077 676 2089 716
rect 2097 676 2109 716
rect 2174 658 2186 716
rect 2210 656 2222 716
rect 2251 676 2263 716
rect 2271 676 2283 716
rect 2291 688 2303 716
rect 2311 676 2323 716
rect 2337 676 2349 716
rect 2357 688 2369 716
rect 2377 676 2389 716
rect 2397 676 2409 716
rect 2438 656 2450 716
rect 2474 658 2486 716
rect 2538 656 2550 716
rect 2574 658 2586 716
rect 2651 696 2663 716
rect 2671 696 2683 716
rect 2698 656 2710 716
rect 2734 658 2746 716
rect 2801 676 2813 716
rect 2821 696 2833 716
rect 2853 696 2865 716
rect 2883 696 2895 716
rect 2905 696 2917 716
rect 2931 696 2943 716
rect 2959 696 2971 716
rect 2989 696 3001 716
rect 3011 676 3023 716
rect 3037 676 3049 716
rect 3057 688 3069 716
rect 3077 676 3089 716
rect 3097 676 3109 716
rect 3137 696 3149 716
rect 3157 696 3169 716
rect 3197 696 3209 716
rect 3217 696 3229 716
rect 3258 656 3270 716
rect 3294 658 3306 716
rect 3371 696 3383 716
rect 3391 696 3403 716
rect 3439 676 3451 716
rect 3469 676 3481 716
rect 3511 676 3523 716
rect 3531 676 3543 716
rect 3551 688 3563 716
rect 3571 676 3583 716
rect 3601 676 3613 716
rect 3621 696 3633 716
rect 3653 696 3665 716
rect 3683 696 3695 716
rect 3705 696 3717 716
rect 3731 696 3743 716
rect 3759 696 3771 716
rect 3789 696 3801 716
rect 3811 676 3823 716
rect 3837 676 3849 716
rect 3857 688 3869 716
rect 3877 676 3889 716
rect 3897 676 3909 716
rect 3959 676 3971 716
rect 3989 676 4001 716
rect 4017 676 4029 716
rect 4039 696 4051 716
rect 4069 696 4081 716
rect 4097 696 4109 716
rect 4123 696 4135 716
rect 4145 696 4157 716
rect 4175 696 4187 716
rect 4207 696 4219 716
rect 4227 676 4239 716
rect 4259 676 4271 716
rect 4289 676 4301 716
rect 4339 676 4351 716
rect 4369 676 4381 716
rect 4431 676 4443 716
rect 4451 676 4463 716
rect 4471 688 4483 716
rect 4491 676 4503 716
rect 4521 676 4533 716
rect 4541 696 4553 716
rect 4573 696 4585 716
rect 4603 696 4615 716
rect 4625 696 4637 716
rect 4651 696 4663 716
rect 4679 696 4691 716
rect 4709 696 4721 716
rect 4731 676 4743 716
rect 19 264 31 304
rect 49 264 61 304
rect 99 264 111 304
rect 129 264 141 304
rect 199 264 211 304
rect 229 264 241 304
rect 279 264 291 304
rect 309 264 321 304
rect 361 264 373 304
rect 381 264 393 304
rect 411 264 423 304
rect 459 264 471 304
rect 489 264 501 304
rect 554 264 566 322
rect 590 264 602 324
rect 652 264 664 304
rect 680 264 692 304
rect 708 264 720 304
rect 751 264 763 284
rect 771 264 783 284
rect 791 264 803 284
rect 839 264 851 304
rect 869 264 881 304
rect 899 264 911 304
rect 929 264 941 304
rect 999 264 1011 304
rect 1029 264 1041 304
rect 1079 264 1091 304
rect 1109 264 1121 304
rect 1172 264 1184 304
rect 1200 264 1212 304
rect 1228 264 1240 304
rect 1257 264 1269 304
rect 1277 264 1289 292
rect 1297 264 1309 304
rect 1317 264 1329 304
rect 1371 264 1383 284
rect 1391 264 1403 284
rect 1411 264 1423 284
rect 1437 264 1449 304
rect 1457 264 1469 292
rect 1477 264 1489 304
rect 1497 264 1509 304
rect 1537 264 1549 284
rect 1557 264 1569 284
rect 1618 264 1630 284
rect 1640 264 1652 304
rect 1668 264 1680 304
rect 1697 264 1709 284
rect 1717 264 1729 284
rect 1758 264 1770 324
rect 1794 264 1806 322
rect 1860 264 1872 304
rect 1888 264 1900 304
rect 1910 264 1922 284
rect 1959 264 1971 304
rect 1989 264 2001 304
rect 2039 264 2051 304
rect 2069 264 2081 304
rect 2119 264 2131 304
rect 2149 264 2161 304
rect 2211 264 2223 284
rect 2231 264 2243 284
rect 2251 264 2263 284
rect 2299 264 2311 304
rect 2329 264 2341 304
rect 2357 264 2369 284
rect 2377 264 2389 284
rect 2397 264 2409 284
rect 2438 264 2450 324
rect 2474 264 2486 322
rect 2551 264 2563 284
rect 2571 264 2583 284
rect 2634 264 2646 322
rect 2670 264 2682 324
rect 2700 264 2712 304
rect 2728 264 2740 304
rect 2750 264 2762 284
rect 2797 264 2809 284
rect 2817 264 2829 284
rect 2837 264 2849 284
rect 2899 264 2911 304
rect 2929 264 2941 304
rect 2971 264 2983 304
rect 2991 264 3003 304
rect 3011 264 3023 292
rect 3031 264 3043 304
rect 3071 264 3083 304
rect 3091 264 3103 304
rect 3111 264 3123 292
rect 3131 264 3143 304
rect 3171 264 3183 284
rect 3191 264 3203 284
rect 3211 264 3223 284
rect 3251 264 3263 284
rect 3271 264 3283 284
rect 3311 264 3323 304
rect 3331 264 3343 304
rect 3351 264 3363 292
rect 3371 264 3383 304
rect 3418 264 3430 284
rect 3440 264 3452 304
rect 3468 264 3480 304
rect 3511 264 3523 284
rect 3531 264 3543 284
rect 3551 264 3563 284
rect 3577 264 3589 284
rect 3597 264 3609 284
rect 3617 264 3629 284
rect 3637 264 3649 304
rect 3679 264 3691 304
rect 3709 264 3721 304
rect 3759 264 3771 304
rect 3789 264 3801 304
rect 3851 264 3863 304
rect 3871 264 3883 304
rect 3891 264 3903 292
rect 3911 264 3923 304
rect 3951 264 3963 284
rect 3971 264 3983 284
rect 4011 264 4023 284
rect 4031 264 4043 284
rect 4057 264 4069 304
rect 4079 264 4091 284
rect 4109 264 4121 284
rect 4137 264 4149 284
rect 4163 264 4175 284
rect 4185 264 4197 284
rect 4215 264 4227 284
rect 4247 264 4259 284
rect 4267 264 4279 304
rect 4319 264 4331 304
rect 4349 264 4361 304
rect 4391 264 4403 304
rect 4411 264 4423 304
rect 4431 264 4443 292
rect 4451 264 4463 304
rect 4491 264 4503 284
rect 4511 264 4523 284
rect 4537 264 4549 304
rect 4559 264 4571 284
rect 4589 264 4601 284
rect 4617 264 4629 284
rect 4643 264 4655 284
rect 4665 264 4677 284
rect 4695 264 4707 284
rect 4727 264 4739 284
rect 4747 264 4759 304
rect 54 178 66 236
rect 90 176 102 236
rect 120 196 132 236
rect 148 196 160 236
rect 170 216 182 236
rect 231 196 243 236
rect 251 196 263 236
rect 271 208 283 236
rect 291 196 303 236
rect 317 196 329 236
rect 337 208 349 236
rect 357 196 369 236
rect 377 196 389 236
rect 454 178 466 236
rect 490 176 502 236
rect 518 176 530 236
rect 554 178 566 236
rect 620 196 632 236
rect 648 196 660 236
rect 670 216 682 236
rect 738 216 750 236
rect 760 196 772 236
rect 788 196 800 236
rect 817 216 829 236
rect 837 216 849 236
rect 891 196 903 236
rect 911 196 923 236
rect 931 208 943 236
rect 951 196 963 236
rect 991 216 1003 236
rect 1011 216 1023 236
rect 1037 196 1049 236
rect 1057 208 1069 236
rect 1077 196 1089 236
rect 1097 196 1109 236
rect 1137 196 1149 236
rect 1157 208 1169 236
rect 1177 196 1189 236
rect 1197 196 1209 236
rect 1238 176 1250 236
rect 1274 178 1286 236
rect 1338 176 1350 236
rect 1374 178 1386 236
rect 1458 216 1470 236
rect 1480 196 1492 236
rect 1508 196 1520 236
rect 1538 176 1550 236
rect 1574 178 1586 236
rect 1658 216 1670 236
rect 1680 196 1692 236
rect 1708 196 1720 236
rect 1738 176 1750 236
rect 1774 178 1786 236
rect 1839 196 1851 236
rect 1869 196 1881 236
rect 1917 216 1929 236
rect 1939 196 1951 236
rect 1959 196 1971 236
rect 2021 196 2033 236
rect 2041 196 2053 236
rect 2071 196 2083 236
rect 2097 216 2109 236
rect 2119 196 2131 236
rect 2139 196 2151 236
rect 2178 176 2190 236
rect 2214 178 2226 236
rect 2280 196 2292 236
rect 2308 196 2320 236
rect 2336 196 2348 236
rect 2397 196 2409 236
rect 2417 208 2429 236
rect 2437 196 2449 236
rect 2457 196 2469 236
rect 2518 216 2530 236
rect 2540 196 2552 236
rect 2568 196 2580 236
rect 2597 196 2609 236
rect 2617 208 2629 236
rect 2637 196 2649 236
rect 2657 196 2669 236
rect 2697 216 2709 236
rect 2717 216 2729 236
rect 2758 176 2770 236
rect 2794 178 2806 236
rect 2857 216 2869 236
rect 2877 216 2889 236
rect 2921 196 2933 236
rect 2941 216 2953 236
rect 2973 216 2985 236
rect 3003 216 3015 236
rect 3025 216 3037 236
rect 3051 216 3063 236
rect 3079 216 3091 236
rect 3109 216 3121 236
rect 3131 196 3143 236
rect 3157 216 3169 236
rect 3177 216 3189 236
rect 3231 216 3243 236
rect 3251 216 3263 236
rect 3281 196 3293 236
rect 3301 216 3313 236
rect 3333 216 3345 236
rect 3363 216 3375 236
rect 3385 216 3397 236
rect 3411 216 3423 236
rect 3439 216 3451 236
rect 3469 216 3481 236
rect 3491 196 3503 236
rect 3531 216 3543 236
rect 3551 216 3563 236
rect 3571 216 3583 236
rect 3597 196 3609 236
rect 3619 216 3631 236
rect 3649 216 3661 236
rect 3677 216 3689 236
rect 3703 216 3715 236
rect 3725 216 3737 236
rect 3755 216 3767 236
rect 3787 216 3799 236
rect 3807 196 3819 236
rect 3837 216 3849 236
rect 3857 216 3869 236
rect 3897 196 3909 236
rect 3917 208 3929 236
rect 3937 196 3949 236
rect 3957 196 3969 236
rect 3997 216 4009 236
rect 4017 216 4029 236
rect 4037 216 4049 236
rect 4077 216 4089 236
rect 4097 216 4109 236
rect 4117 216 4129 236
rect 4171 216 4183 236
rect 4191 216 4203 236
rect 4211 216 4223 236
rect 4237 196 4249 236
rect 4257 208 4269 236
rect 4277 196 4289 236
rect 4297 196 4309 236
rect 4359 196 4371 236
rect 4389 196 4401 236
rect 4431 216 4443 236
rect 4451 216 4463 236
rect 4477 216 4489 236
rect 4497 216 4509 236
rect 4517 216 4529 236
rect 4559 196 4571 236
rect 4589 196 4601 236
rect 4651 216 4663 236
rect 4671 216 4683 236
rect 4699 196 4711 236
rect 4729 196 4741 236
<< pdcontact >>
rect 31 4344 43 4424
rect 51 4344 63 4424
rect 71 4344 83 4412
rect 91 4344 103 4416
rect 131 4344 143 4384
rect 151 4344 163 4380
rect 171 4344 183 4384
rect 191 4344 203 4384
rect 217 4344 229 4384
rect 237 4344 249 4384
rect 257 4344 269 4380
rect 277 4344 289 4384
rect 331 4344 343 4384
rect 351 4344 363 4380
rect 371 4344 383 4384
rect 391 4344 403 4384
rect 417 4344 429 4416
rect 437 4344 449 4412
rect 457 4344 469 4424
rect 477 4344 489 4424
rect 522 4344 534 4424
rect 550 4344 562 4424
rect 572 4344 584 4384
rect 622 4344 634 4424
rect 650 4344 662 4424
rect 672 4344 684 4384
rect 731 4344 743 4384
rect 751 4344 763 4380
rect 771 4344 783 4384
rect 791 4344 803 4384
rect 817 4344 829 4384
rect 837 4344 849 4384
rect 857 4344 869 4380
rect 877 4344 889 4384
rect 917 4344 929 4384
rect 937 4344 949 4384
rect 957 4344 969 4384
rect 997 4344 1009 4384
rect 1017 4344 1029 4384
rect 1037 4344 1049 4380
rect 1057 4344 1069 4384
rect 1097 4344 1109 4416
rect 1117 4344 1129 4412
rect 1137 4344 1149 4424
rect 1157 4344 1169 4424
rect 1211 4344 1223 4384
rect 1231 4344 1243 4384
rect 1251 4344 1263 4384
rect 1303 4344 1315 4424
rect 1331 4344 1343 4424
rect 1376 4344 1388 4384
rect 1398 4344 1410 4424
rect 1426 4344 1438 4424
rect 1471 4344 1483 4384
rect 1491 4344 1503 4384
rect 1511 4344 1523 4384
rect 1537 4344 1549 4424
rect 1565 4344 1577 4424
rect 1617 4344 1629 4384
rect 1637 4344 1649 4384
rect 1657 4344 1669 4380
rect 1677 4344 1689 4384
rect 1731 4344 1743 4424
rect 1751 4344 1763 4424
rect 1771 4344 1783 4412
rect 1791 4344 1803 4416
rect 1817 4344 1829 4384
rect 1837 4344 1849 4384
rect 1891 4344 1903 4384
rect 1911 4344 1923 4384
rect 1937 4344 1949 4416
rect 1957 4344 1969 4412
rect 1977 4344 1989 4424
rect 1997 4344 2009 4424
rect 2037 4344 2049 4424
rect 2065 4344 2077 4424
rect 2117 4344 2129 4384
rect 2137 4344 2149 4384
rect 2182 4344 2194 4424
rect 2210 4344 2222 4424
rect 2232 4344 2244 4384
rect 2301 4344 2313 4424
rect 2331 4344 2353 4424
rect 2371 4344 2383 4424
rect 2397 4344 2409 4424
rect 2427 4344 2439 4423
rect 2447 4344 2459 4423
rect 2497 4344 2509 4416
rect 2517 4344 2529 4412
rect 2537 4344 2549 4424
rect 2557 4344 2569 4424
rect 2611 4344 2623 4424
rect 2631 4356 2643 4424
rect 2651 4344 2663 4422
rect 2671 4344 2683 4410
rect 2691 4344 2703 4422
rect 2721 4344 2733 4424
rect 2741 4344 2753 4384
rect 2775 4344 2787 4384
rect 2807 4344 2819 4384
rect 2827 4344 2839 4384
rect 2853 4344 2865 4384
rect 2881 4344 2893 4364
rect 2911 4344 2923 4364
rect 2931 4344 2943 4424
rect 2971 4344 2983 4384
rect 2991 4344 3003 4384
rect 3036 4344 3048 4384
rect 3058 4344 3070 4424
rect 3086 4344 3098 4424
rect 3143 4344 3155 4424
rect 3171 4344 3183 4424
rect 3216 4344 3228 4384
rect 3238 4344 3250 4424
rect 3266 4344 3278 4424
rect 3323 4344 3335 4424
rect 3351 4344 3363 4424
rect 3391 4344 3403 4384
rect 3411 4344 3423 4384
rect 3437 4344 3449 4424
rect 3457 4344 3469 4364
rect 3487 4344 3499 4364
rect 3515 4344 3527 4384
rect 3541 4344 3553 4384
rect 3561 4344 3573 4384
rect 3593 4344 3605 4384
rect 3627 4344 3639 4384
rect 3647 4344 3659 4424
rect 3682 4344 3694 4424
rect 3710 4344 3722 4424
rect 3732 4344 3744 4384
rect 3777 4344 3789 4384
rect 3797 4344 3809 4384
rect 3817 4344 3829 4384
rect 3871 4344 3883 4424
rect 3891 4344 3903 4424
rect 3911 4344 3923 4424
rect 3931 4344 3943 4424
rect 3951 4344 3963 4424
rect 3971 4344 3983 4424
rect 3991 4344 4003 4424
rect 4011 4344 4023 4424
rect 4031 4344 4043 4424
rect 4069 4344 4081 4424
rect 4089 4344 4101 4424
rect 4111 4344 4123 4384
rect 4137 4344 4149 4384
rect 4157 4344 4169 4384
rect 4177 4344 4189 4384
rect 4217 4344 4229 4384
rect 4237 4344 4249 4384
rect 4282 4344 4294 4424
rect 4310 4344 4322 4424
rect 4332 4344 4344 4384
rect 4377 4344 4389 4424
rect 4397 4344 4409 4364
rect 4427 4344 4439 4364
rect 4455 4344 4467 4384
rect 4481 4344 4493 4384
rect 4501 4344 4513 4384
rect 4533 4344 4545 4384
rect 4567 4344 4579 4384
rect 4587 4344 4599 4424
rect 4617 4344 4629 4384
rect 4639 4344 4651 4424
rect 4659 4344 4671 4424
rect 4697 4344 4709 4384
rect 4717 4344 4729 4384
rect 4737 4344 4749 4384
rect 31 4276 43 4316
rect 51 4276 63 4316
rect 71 4276 83 4316
rect 97 4244 109 4316
rect 117 4248 129 4316
rect 137 4236 149 4316
rect 157 4236 169 4316
rect 211 4276 223 4316
rect 231 4276 243 4316
rect 251 4276 263 4316
rect 303 4236 315 4316
rect 331 4236 343 4316
rect 376 4276 388 4316
rect 398 4236 410 4316
rect 426 4236 438 4316
rect 462 4236 474 4316
rect 490 4236 502 4316
rect 512 4276 524 4316
rect 571 4276 583 4316
rect 591 4276 603 4316
rect 631 4236 643 4316
rect 651 4236 663 4316
rect 671 4248 683 4316
rect 691 4244 703 4316
rect 731 4276 743 4316
rect 751 4276 763 4316
rect 777 4276 789 4316
rect 797 4276 809 4316
rect 817 4280 829 4316
rect 837 4276 849 4316
rect 891 4236 903 4316
rect 911 4236 923 4304
rect 931 4238 943 4316
rect 951 4250 963 4316
rect 971 4238 983 4316
rect 1011 4276 1023 4316
rect 1031 4280 1043 4316
rect 1051 4276 1063 4316
rect 1071 4276 1083 4316
rect 1097 4276 1109 4316
rect 1117 4276 1129 4316
rect 1137 4280 1149 4316
rect 1157 4276 1169 4316
rect 1211 4276 1223 4316
rect 1231 4276 1243 4316
rect 1251 4276 1263 4316
rect 1291 4276 1303 4316
rect 1311 4280 1323 4316
rect 1331 4276 1343 4316
rect 1351 4276 1363 4316
rect 1391 4276 1403 4316
rect 1411 4276 1423 4316
rect 1431 4276 1443 4316
rect 1457 4276 1469 4316
rect 1477 4276 1489 4316
rect 1497 4280 1509 4316
rect 1517 4276 1529 4316
rect 1583 4236 1595 4316
rect 1611 4236 1623 4316
rect 1663 4236 1675 4316
rect 1691 4236 1703 4316
rect 1722 4236 1734 4316
rect 1750 4236 1762 4316
rect 1772 4276 1784 4316
rect 1831 4276 1843 4316
rect 1851 4276 1863 4316
rect 1871 4276 1883 4316
rect 1897 4276 1909 4316
rect 1917 4276 1929 4316
rect 1957 4276 1969 4316
rect 1977 4276 1989 4316
rect 1997 4280 2009 4316
rect 2017 4276 2029 4316
rect 2057 4276 2069 4316
rect 2077 4276 2089 4316
rect 2097 4280 2109 4316
rect 2117 4276 2129 4316
rect 2161 4236 2173 4316
rect 2181 4276 2193 4316
rect 2215 4276 2227 4316
rect 2247 4276 2259 4316
rect 2267 4276 2279 4316
rect 2293 4276 2305 4316
rect 2321 4296 2333 4316
rect 2351 4296 2363 4316
rect 2371 4236 2383 4316
rect 2397 4276 2409 4316
rect 2419 4236 2431 4316
rect 2439 4236 2451 4316
rect 2491 4276 2503 4316
rect 2511 4276 2523 4316
rect 2563 4236 2575 4316
rect 2591 4236 2603 4316
rect 2617 4236 2629 4316
rect 2637 4296 2649 4316
rect 2667 4296 2679 4316
rect 2695 4276 2707 4316
rect 2721 4276 2733 4316
rect 2741 4276 2753 4316
rect 2773 4276 2785 4316
rect 2807 4276 2819 4316
rect 2827 4236 2839 4316
rect 2857 4276 2869 4316
rect 2877 4276 2889 4316
rect 2943 4236 2955 4316
rect 2971 4236 2983 4316
rect 3002 4236 3014 4316
rect 3030 4236 3042 4316
rect 3052 4276 3064 4316
rect 3097 4276 3109 4316
rect 3117 4276 3129 4316
rect 3137 4276 3149 4316
rect 3191 4276 3203 4316
rect 3211 4276 3223 4316
rect 3231 4276 3243 4316
rect 3271 4276 3283 4316
rect 3291 4276 3303 4316
rect 3311 4276 3323 4316
rect 3337 4236 3349 4316
rect 3365 4236 3377 4316
rect 3421 4236 3433 4316
rect 3441 4276 3453 4316
rect 3475 4276 3487 4316
rect 3507 4276 3519 4316
rect 3527 4276 3539 4316
rect 3553 4276 3565 4316
rect 3581 4296 3593 4316
rect 3611 4296 3623 4316
rect 3631 4236 3643 4316
rect 3671 4276 3683 4316
rect 3691 4276 3703 4316
rect 3711 4276 3723 4316
rect 3737 4236 3749 4316
rect 3765 4236 3777 4316
rect 3817 4236 3829 4316
rect 3837 4296 3849 4316
rect 3867 4296 3879 4316
rect 3895 4276 3907 4316
rect 3921 4276 3933 4316
rect 3941 4276 3953 4316
rect 3973 4276 3985 4316
rect 4007 4276 4019 4316
rect 4027 4236 4039 4316
rect 4057 4236 4069 4316
rect 4085 4236 4097 4316
rect 4151 4236 4163 4316
rect 4171 4236 4183 4316
rect 4191 4248 4203 4316
rect 4211 4244 4223 4316
rect 4237 4276 4249 4316
rect 4259 4236 4271 4316
rect 4279 4236 4291 4316
rect 4343 4236 4355 4316
rect 4371 4236 4383 4316
rect 4411 4236 4423 4316
rect 4431 4236 4443 4316
rect 4451 4248 4463 4316
rect 4471 4244 4483 4316
rect 4497 4236 4509 4316
rect 4517 4296 4529 4316
rect 4547 4296 4559 4316
rect 4575 4276 4587 4316
rect 4601 4276 4613 4316
rect 4621 4276 4633 4316
rect 4653 4276 4665 4316
rect 4687 4276 4699 4316
rect 4707 4236 4719 4316
rect 31 3864 43 3904
rect 51 3864 63 3904
rect 71 3864 83 3904
rect 97 3864 109 3904
rect 117 3864 129 3904
rect 137 3864 149 3904
rect 191 3864 203 3904
rect 211 3864 223 3904
rect 231 3864 243 3904
rect 276 3864 288 3904
rect 298 3864 310 3944
rect 326 3864 338 3944
rect 357 3864 369 3936
rect 377 3864 389 3932
rect 397 3864 409 3944
rect 417 3864 429 3944
rect 483 3864 495 3944
rect 511 3864 523 3944
rect 537 3864 549 3904
rect 557 3864 569 3904
rect 577 3864 589 3904
rect 622 3864 634 3944
rect 650 3864 662 3944
rect 672 3864 684 3904
rect 731 3864 743 3904
rect 751 3864 763 3900
rect 771 3864 783 3904
rect 791 3864 803 3904
rect 817 3864 829 3904
rect 837 3864 849 3904
rect 857 3864 869 3900
rect 877 3864 889 3904
rect 936 3864 948 3904
rect 958 3864 970 3944
rect 986 3864 998 3944
rect 1022 3864 1034 3944
rect 1050 3864 1062 3944
rect 1072 3864 1084 3904
rect 1131 3864 1143 3904
rect 1151 3864 1163 3904
rect 1191 3864 1203 3904
rect 1211 3864 1223 3900
rect 1231 3864 1243 3904
rect 1251 3864 1263 3904
rect 1277 3864 1289 3904
rect 1297 3864 1309 3904
rect 1337 3864 1349 3904
rect 1357 3864 1369 3904
rect 1377 3864 1389 3900
rect 1397 3864 1409 3904
rect 1437 3864 1449 3904
rect 1457 3864 1469 3904
rect 1477 3864 1489 3900
rect 1497 3864 1509 3904
rect 1537 3864 1549 3904
rect 1557 3864 1569 3904
rect 1577 3864 1589 3904
rect 1643 3864 1655 3944
rect 1671 3864 1683 3944
rect 1707 3864 1719 3944
rect 1727 3864 1739 3944
rect 1751 3864 1763 3904
rect 1771 3864 1783 3904
rect 1816 3864 1828 3904
rect 1838 3864 1850 3944
rect 1866 3864 1878 3944
rect 1897 3864 1909 3944
rect 1925 3864 1937 3944
rect 1991 3864 2003 3904
rect 2011 3864 2023 3904
rect 2042 3864 2054 3944
rect 2070 3864 2082 3944
rect 2092 3864 2104 3904
rect 2137 3864 2149 3904
rect 2157 3864 2169 3904
rect 2197 3864 2209 3904
rect 2217 3864 2229 3904
rect 2237 3864 2249 3904
rect 2277 3864 2289 3904
rect 2297 3864 2309 3904
rect 2317 3864 2329 3900
rect 2337 3864 2349 3904
rect 2377 3864 2389 3904
rect 2399 3864 2411 3944
rect 2419 3864 2431 3944
rect 2457 3864 2469 3944
rect 2477 3864 2489 3944
rect 2497 3864 2509 3944
rect 2517 3864 2529 3944
rect 2537 3864 2549 3944
rect 2557 3864 2569 3944
rect 2577 3864 2589 3944
rect 2597 3864 2609 3944
rect 2617 3864 2629 3944
rect 2661 3864 2673 3944
rect 2681 3864 2693 3904
rect 2715 3864 2727 3904
rect 2747 3864 2759 3904
rect 2767 3864 2779 3904
rect 2793 3864 2805 3904
rect 2821 3864 2833 3884
rect 2851 3864 2863 3884
rect 2871 3864 2883 3944
rect 2897 3864 2909 3904
rect 2917 3864 2929 3904
rect 2962 3864 2974 3944
rect 2990 3864 3002 3944
rect 3012 3864 3024 3904
rect 3057 3864 3069 3944
rect 3085 3864 3097 3944
rect 3137 3864 3149 3904
rect 3157 3864 3169 3904
rect 3177 3864 3189 3904
rect 3231 3864 3243 3944
rect 3251 3864 3263 3944
rect 3271 3864 3283 3932
rect 3291 3864 3303 3936
rect 3317 3864 3329 3904
rect 3337 3864 3349 3904
rect 3361 3864 3373 3944
rect 3381 3864 3393 3944
rect 3443 3864 3455 3944
rect 3471 3864 3483 3944
rect 3511 3864 3523 3904
rect 3531 3864 3543 3904
rect 3557 3864 3569 3944
rect 3577 3864 3589 3884
rect 3607 3864 3619 3884
rect 3635 3864 3647 3904
rect 3661 3864 3673 3904
rect 3681 3864 3693 3904
rect 3713 3864 3725 3904
rect 3747 3864 3759 3904
rect 3767 3864 3779 3944
rect 3811 3864 3823 3944
rect 3831 3864 3843 3944
rect 3851 3864 3863 3932
rect 3871 3864 3883 3936
rect 3897 3864 3909 3944
rect 3925 3864 3937 3944
rect 4003 3864 4015 3944
rect 4031 3864 4043 3944
rect 4057 3864 4069 3904
rect 4077 3864 4089 3904
rect 4101 3864 4113 3944
rect 4121 3864 4133 3944
rect 4162 3864 4174 3944
rect 4190 3864 4202 3944
rect 4212 3864 4224 3904
rect 4276 3864 4288 3904
rect 4298 3864 4310 3944
rect 4326 3864 4338 3944
rect 4371 3864 4383 3904
rect 4391 3864 4403 3904
rect 4417 3864 4429 3944
rect 4437 3864 4449 3884
rect 4467 3864 4479 3884
rect 4495 3864 4507 3904
rect 4521 3864 4533 3904
rect 4541 3864 4553 3904
rect 4573 3864 4585 3904
rect 4607 3864 4619 3904
rect 4627 3864 4639 3944
rect 4657 3864 4669 3904
rect 4677 3864 4689 3904
rect 43 3756 55 3836
rect 71 3756 83 3836
rect 102 3756 114 3836
rect 130 3756 142 3836
rect 152 3796 164 3836
rect 211 3796 223 3836
rect 231 3796 243 3836
rect 271 3756 283 3836
rect 291 3756 303 3836
rect 311 3768 323 3836
rect 331 3764 343 3836
rect 367 3756 379 3836
rect 387 3756 399 3836
rect 411 3796 423 3836
rect 431 3796 443 3836
rect 471 3796 483 3836
rect 491 3796 503 3836
rect 511 3796 523 3836
rect 551 3796 563 3836
rect 571 3796 583 3836
rect 591 3796 603 3836
rect 617 3796 629 3836
rect 637 3796 649 3836
rect 682 3756 694 3836
rect 710 3756 722 3836
rect 732 3796 744 3836
rect 777 3796 789 3836
rect 797 3796 809 3836
rect 817 3796 829 3836
rect 871 3796 883 3836
rect 891 3800 903 3836
rect 911 3796 923 3836
rect 931 3796 943 3836
rect 957 3764 969 3836
rect 977 3768 989 3836
rect 997 3756 1009 3836
rect 1017 3756 1029 3836
rect 1057 3796 1069 3836
rect 1077 3796 1089 3836
rect 1097 3800 1109 3836
rect 1117 3796 1129 3836
rect 1157 3764 1169 3836
rect 1177 3768 1189 3836
rect 1197 3756 1209 3836
rect 1217 3756 1229 3836
rect 1257 3796 1269 3836
rect 1277 3796 1289 3836
rect 1331 3796 1343 3836
rect 1351 3800 1363 3836
rect 1371 3796 1383 3836
rect 1391 3796 1403 3836
rect 1431 3796 1443 3836
rect 1451 3796 1463 3836
rect 1496 3796 1508 3836
rect 1518 3756 1530 3836
rect 1546 3756 1558 3836
rect 1591 3796 1603 3836
rect 1611 3796 1623 3836
rect 1637 3764 1649 3836
rect 1657 3768 1669 3836
rect 1677 3756 1689 3836
rect 1697 3756 1709 3836
rect 1737 3756 1749 3836
rect 1765 3756 1777 3836
rect 1831 3756 1843 3836
rect 1851 3756 1863 3836
rect 1871 3768 1883 3836
rect 1891 3764 1903 3836
rect 1931 3796 1943 3836
rect 1951 3796 1963 3836
rect 1971 3796 1983 3836
rect 1997 3756 2009 3836
rect 2027 3757 2039 3836
rect 2047 3757 2059 3836
rect 2097 3796 2109 3836
rect 2119 3756 2131 3836
rect 2139 3756 2151 3836
rect 2191 3756 2203 3836
rect 2211 3756 2223 3836
rect 2231 3756 2243 3836
rect 2251 3756 2263 3836
rect 2271 3756 2283 3836
rect 2291 3756 2303 3836
rect 2311 3756 2323 3836
rect 2331 3756 2343 3836
rect 2351 3756 2363 3836
rect 2381 3756 2393 3836
rect 2401 3796 2413 3836
rect 2435 3796 2447 3836
rect 2467 3796 2479 3836
rect 2487 3796 2499 3836
rect 2513 3796 2525 3836
rect 2541 3816 2553 3836
rect 2571 3816 2583 3836
rect 2591 3756 2603 3836
rect 2636 3796 2648 3836
rect 2658 3756 2670 3836
rect 2686 3756 2698 3836
rect 2731 3796 2743 3836
rect 2751 3796 2763 3836
rect 2803 3756 2815 3836
rect 2831 3756 2843 3836
rect 2883 3756 2895 3836
rect 2911 3756 2923 3836
rect 2963 3756 2975 3836
rect 2991 3756 3003 3836
rect 3017 3796 3029 3836
rect 3037 3796 3049 3836
rect 3091 3796 3103 3836
rect 3111 3796 3123 3836
rect 3142 3756 3154 3836
rect 3170 3756 3182 3836
rect 3192 3796 3204 3836
rect 3251 3756 3263 3836
rect 3271 3756 3283 3836
rect 3291 3768 3303 3836
rect 3311 3764 3323 3836
rect 3337 3764 3349 3836
rect 3357 3768 3369 3836
rect 3377 3756 3389 3836
rect 3397 3756 3409 3836
rect 3437 3796 3449 3836
rect 3457 3796 3469 3836
rect 3497 3796 3509 3836
rect 3517 3796 3529 3836
rect 3541 3756 3553 3836
rect 3561 3756 3573 3836
rect 3602 3756 3614 3836
rect 3630 3756 3642 3836
rect 3652 3796 3664 3836
rect 3702 3756 3714 3836
rect 3730 3756 3742 3836
rect 3752 3796 3764 3836
rect 3801 3756 3813 3836
rect 3821 3796 3833 3836
rect 3855 3796 3867 3836
rect 3887 3796 3899 3836
rect 3907 3796 3919 3836
rect 3933 3796 3945 3836
rect 3961 3816 3973 3836
rect 3991 3816 4003 3836
rect 4011 3756 4023 3836
rect 4037 3796 4049 3836
rect 4059 3756 4071 3836
rect 4079 3756 4091 3836
rect 4143 3756 4155 3836
rect 4171 3756 4183 3836
rect 4197 3764 4209 3836
rect 4217 3768 4229 3836
rect 4237 3756 4249 3836
rect 4257 3756 4269 3836
rect 4297 3756 4309 3836
rect 4317 3816 4329 3836
rect 4347 3816 4359 3836
rect 4375 3796 4387 3836
rect 4401 3796 4413 3836
rect 4421 3796 4433 3836
rect 4453 3796 4465 3836
rect 4487 3796 4499 3836
rect 4507 3756 4519 3836
rect 4537 3796 4549 3836
rect 4559 3756 4571 3836
rect 4579 3756 4591 3836
rect 4631 3796 4643 3836
rect 4651 3796 4663 3836
rect 4677 3796 4689 3836
rect 4697 3796 4709 3836
rect 31 3384 43 3424
rect 51 3384 63 3424
rect 71 3384 83 3424
rect 101 3384 113 3464
rect 121 3384 133 3424
rect 155 3384 167 3424
rect 187 3384 199 3424
rect 207 3384 219 3424
rect 233 3384 245 3424
rect 261 3384 273 3404
rect 291 3384 303 3404
rect 311 3384 323 3464
rect 351 3384 363 3424
rect 371 3384 383 3424
rect 411 3384 423 3424
rect 431 3384 443 3424
rect 451 3384 463 3424
rect 496 3384 508 3424
rect 518 3384 530 3464
rect 546 3384 558 3464
rect 596 3384 608 3424
rect 618 3384 630 3464
rect 646 3384 658 3464
rect 677 3384 689 3424
rect 697 3384 709 3424
rect 717 3384 729 3424
rect 757 3384 769 3464
rect 787 3384 809 3464
rect 827 3384 839 3464
rect 877 3384 889 3424
rect 897 3384 909 3424
rect 951 3384 963 3424
rect 971 3384 983 3420
rect 991 3384 1003 3424
rect 1011 3384 1023 3424
rect 1037 3384 1049 3456
rect 1057 3384 1069 3452
rect 1077 3384 1089 3464
rect 1097 3384 1109 3464
rect 1137 3384 1149 3464
rect 1165 3384 1177 3464
rect 1217 3384 1229 3424
rect 1237 3384 1249 3424
rect 1257 3384 1269 3424
rect 1297 3384 1309 3424
rect 1317 3384 1329 3424
rect 1337 3384 1349 3424
rect 1382 3384 1394 3464
rect 1410 3384 1422 3464
rect 1432 3384 1444 3424
rect 1481 3384 1493 3464
rect 1501 3384 1513 3424
rect 1535 3384 1547 3424
rect 1567 3384 1579 3424
rect 1587 3384 1599 3424
rect 1613 3384 1625 3424
rect 1641 3384 1653 3404
rect 1671 3384 1683 3404
rect 1691 3384 1703 3464
rect 1731 3384 1743 3424
rect 1751 3384 1763 3424
rect 1771 3384 1783 3424
rect 1802 3384 1814 3464
rect 1830 3384 1842 3464
rect 1852 3384 1864 3424
rect 1897 3384 1909 3464
rect 1917 3384 1929 3464
rect 1971 3384 1983 3424
rect 1991 3384 2003 3424
rect 2011 3384 2023 3424
rect 2047 3384 2059 3464
rect 2067 3384 2079 3464
rect 2091 3384 2103 3424
rect 2111 3384 2123 3424
rect 2137 3384 2149 3424
rect 2157 3384 2169 3424
rect 2177 3384 2189 3424
rect 2217 3384 2229 3424
rect 2237 3384 2249 3424
rect 2257 3384 2269 3420
rect 2277 3384 2289 3424
rect 2317 3384 2329 3424
rect 2337 3384 2349 3424
rect 2377 3384 2389 3424
rect 2397 3384 2409 3424
rect 2437 3384 2449 3464
rect 2457 3384 2469 3404
rect 2487 3384 2499 3404
rect 2515 3384 2527 3424
rect 2541 3384 2553 3424
rect 2561 3384 2573 3424
rect 2593 3384 2605 3424
rect 2627 3384 2639 3424
rect 2647 3384 2659 3464
rect 2682 3384 2694 3464
rect 2710 3384 2722 3464
rect 2732 3384 2744 3424
rect 2777 3384 2789 3424
rect 2799 3384 2811 3464
rect 2819 3384 2831 3464
rect 2857 3384 2869 3424
rect 2877 3384 2889 3424
rect 2897 3384 2909 3424
rect 2937 3384 2949 3464
rect 2957 3384 2969 3404
rect 2987 3384 2999 3404
rect 3015 3384 3027 3424
rect 3041 3384 3053 3424
rect 3061 3384 3073 3424
rect 3093 3384 3105 3424
rect 3127 3384 3139 3424
rect 3147 3384 3159 3464
rect 3196 3384 3208 3424
rect 3218 3384 3230 3464
rect 3246 3384 3258 3464
rect 3291 3384 3303 3424
rect 3311 3384 3323 3424
rect 3337 3384 3349 3464
rect 3365 3384 3377 3464
rect 3417 3384 3429 3424
rect 3437 3384 3449 3424
rect 3503 3384 3515 3464
rect 3531 3384 3543 3464
rect 3557 3384 3569 3456
rect 3577 3384 3589 3452
rect 3597 3384 3609 3464
rect 3617 3384 3629 3464
rect 3657 3384 3669 3464
rect 3687 3384 3699 3463
rect 3707 3384 3719 3463
rect 3771 3384 3783 3464
rect 3791 3396 3803 3464
rect 3811 3384 3823 3462
rect 3831 3384 3843 3450
rect 3851 3384 3863 3462
rect 3891 3384 3903 3424
rect 3911 3384 3923 3424
rect 3931 3384 3943 3424
rect 3957 3384 3969 3464
rect 3977 3384 3989 3404
rect 4007 3384 4019 3404
rect 4035 3384 4047 3424
rect 4061 3384 4073 3424
rect 4081 3384 4093 3424
rect 4113 3384 4125 3424
rect 4147 3384 4159 3424
rect 4167 3384 4179 3464
rect 4197 3384 4209 3464
rect 4217 3384 4229 3404
rect 4247 3384 4259 3404
rect 4275 3384 4287 3424
rect 4301 3384 4313 3424
rect 4321 3384 4333 3424
rect 4353 3384 4365 3424
rect 4387 3384 4399 3424
rect 4407 3384 4419 3464
rect 4451 3384 4463 3464
rect 4471 3384 4483 3464
rect 4491 3384 4503 3464
rect 4511 3384 4523 3464
rect 4531 3384 4543 3464
rect 4551 3384 4563 3464
rect 4571 3384 4583 3464
rect 4591 3384 4603 3464
rect 4611 3384 4623 3464
rect 4642 3384 4654 3464
rect 4670 3384 4682 3464
rect 4692 3384 4704 3424
rect 21 3276 33 3356
rect 41 3316 53 3356
rect 75 3316 87 3356
rect 107 3316 119 3356
rect 127 3316 139 3356
rect 153 3316 165 3356
rect 181 3336 193 3356
rect 211 3336 223 3356
rect 231 3276 243 3356
rect 271 3276 283 3356
rect 291 3276 303 3344
rect 311 3278 323 3356
rect 331 3290 343 3356
rect 351 3278 363 3356
rect 391 3316 403 3356
rect 411 3316 423 3356
rect 431 3316 443 3356
rect 457 3276 469 3356
rect 477 3336 489 3356
rect 507 3336 519 3356
rect 535 3316 547 3356
rect 561 3316 573 3356
rect 581 3316 593 3356
rect 613 3316 625 3356
rect 647 3316 659 3356
rect 667 3276 679 3356
rect 716 3316 728 3356
rect 738 3276 750 3356
rect 766 3276 778 3356
rect 811 3276 823 3356
rect 831 3276 843 3344
rect 851 3278 863 3356
rect 871 3290 883 3356
rect 891 3278 903 3356
rect 917 3316 929 3356
rect 937 3316 949 3356
rect 957 3316 969 3356
rect 1011 3316 1023 3356
rect 1031 3320 1043 3356
rect 1051 3316 1063 3356
rect 1071 3316 1083 3356
rect 1107 3276 1119 3356
rect 1127 3276 1139 3356
rect 1151 3316 1163 3356
rect 1171 3316 1183 3356
rect 1197 3316 1209 3356
rect 1217 3316 1229 3356
rect 1237 3320 1249 3356
rect 1257 3316 1269 3356
rect 1302 3276 1314 3356
rect 1330 3276 1342 3356
rect 1352 3316 1364 3356
rect 1397 3316 1409 3356
rect 1417 3316 1429 3356
rect 1437 3316 1449 3356
rect 1501 3277 1513 3356
rect 1521 3277 1533 3356
rect 1551 3276 1563 3356
rect 1591 3316 1603 3356
rect 1611 3316 1623 3356
rect 1631 3316 1643 3356
rect 1662 3276 1674 3356
rect 1690 3276 1702 3356
rect 1712 3316 1724 3356
rect 1776 3316 1788 3356
rect 1798 3276 1810 3356
rect 1826 3276 1838 3356
rect 1857 3316 1869 3356
rect 1877 3316 1889 3356
rect 1897 3316 1909 3356
rect 1942 3276 1954 3356
rect 1970 3276 1982 3356
rect 1992 3316 2004 3356
rect 2056 3316 2068 3356
rect 2078 3276 2090 3356
rect 2106 3276 2118 3356
rect 2137 3316 2149 3356
rect 2157 3316 2169 3356
rect 2202 3276 2214 3356
rect 2230 3276 2242 3356
rect 2252 3316 2264 3356
rect 2311 3316 2323 3356
rect 2331 3316 2343 3356
rect 2357 3316 2369 3356
rect 2377 3316 2389 3356
rect 2397 3316 2409 3356
rect 2437 3276 2449 3356
rect 2457 3336 2469 3356
rect 2487 3336 2499 3356
rect 2515 3316 2527 3356
rect 2541 3316 2553 3356
rect 2561 3316 2573 3356
rect 2593 3316 2605 3356
rect 2627 3316 2639 3356
rect 2647 3276 2659 3356
rect 2677 3316 2689 3356
rect 2699 3276 2711 3356
rect 2719 3276 2731 3356
rect 2757 3276 2769 3356
rect 2777 3336 2789 3356
rect 2807 3336 2819 3356
rect 2835 3316 2847 3356
rect 2861 3316 2873 3356
rect 2881 3316 2893 3356
rect 2913 3316 2925 3356
rect 2947 3316 2959 3356
rect 2967 3276 2979 3356
rect 3016 3316 3028 3356
rect 3038 3276 3050 3356
rect 3066 3276 3078 3356
rect 3116 3316 3128 3356
rect 3138 3276 3150 3356
rect 3166 3276 3178 3356
rect 3202 3276 3214 3356
rect 3230 3276 3242 3356
rect 3252 3316 3264 3356
rect 3316 3316 3328 3356
rect 3338 3276 3350 3356
rect 3366 3276 3378 3356
rect 3402 3276 3414 3356
rect 3430 3276 3442 3356
rect 3452 3316 3464 3356
rect 3497 3316 3509 3356
rect 3517 3316 3529 3356
rect 3537 3316 3549 3356
rect 3577 3316 3589 3356
rect 3597 3316 3609 3356
rect 3617 3316 3629 3356
rect 3657 3316 3669 3356
rect 3677 3316 3689 3356
rect 3697 3316 3709 3356
rect 3737 3316 3749 3356
rect 3757 3316 3769 3356
rect 3777 3316 3789 3356
rect 3817 3316 3829 3356
rect 3839 3276 3851 3356
rect 3859 3276 3871 3356
rect 3911 3316 3923 3356
rect 3931 3316 3943 3356
rect 3951 3316 3963 3356
rect 4003 3276 4015 3356
rect 4031 3276 4043 3356
rect 4057 3316 4069 3356
rect 4079 3276 4091 3356
rect 4099 3276 4111 3356
rect 4151 3316 4163 3356
rect 4171 3316 4183 3356
rect 4216 3316 4228 3356
rect 4238 3276 4250 3356
rect 4266 3276 4278 3356
rect 4311 3316 4323 3356
rect 4331 3316 4343 3356
rect 4362 3276 4374 3356
rect 4390 3276 4402 3356
rect 4412 3316 4424 3356
rect 4471 3316 4483 3356
rect 4491 3316 4503 3356
rect 4511 3316 4523 3356
rect 4541 3276 4553 3356
rect 4561 3316 4573 3356
rect 4595 3316 4607 3356
rect 4627 3316 4639 3356
rect 4647 3316 4659 3356
rect 4673 3316 4685 3356
rect 4701 3336 4713 3356
rect 4731 3336 4743 3356
rect 4751 3276 4763 3356
rect 31 2904 43 2984
rect 51 2916 63 2984
rect 71 2904 83 2982
rect 91 2904 103 2970
rect 111 2904 123 2982
rect 147 2904 159 2984
rect 167 2904 179 2984
rect 191 2904 203 2944
rect 211 2904 223 2944
rect 237 2904 249 2984
rect 257 2904 269 2924
rect 287 2904 299 2924
rect 315 2904 327 2944
rect 341 2904 353 2944
rect 361 2904 373 2944
rect 393 2904 405 2944
rect 427 2904 439 2944
rect 447 2904 459 2984
rect 482 2904 494 2984
rect 510 2904 522 2984
rect 532 2904 544 2944
rect 577 2904 589 2944
rect 597 2904 609 2944
rect 617 2904 629 2944
rect 671 2904 683 2944
rect 691 2904 703 2944
rect 711 2904 723 2944
rect 763 2904 775 2984
rect 791 2904 803 2984
rect 817 2904 829 2944
rect 837 2904 849 2944
rect 857 2904 869 2944
rect 916 2904 928 2944
rect 938 2904 950 2984
rect 966 2904 978 2984
rect 1016 2904 1028 2944
rect 1038 2904 1050 2984
rect 1066 2904 1078 2984
rect 1123 2904 1135 2984
rect 1151 2904 1163 2984
rect 1196 2904 1208 2944
rect 1218 2904 1230 2984
rect 1246 2904 1258 2984
rect 1277 2904 1289 2944
rect 1297 2904 1309 2944
rect 1317 2904 1329 2944
rect 1371 2904 1383 2984
rect 1391 2904 1403 2984
rect 1417 2904 1429 2944
rect 1437 2904 1449 2944
rect 1457 2904 1469 2944
rect 1497 2904 1509 2944
rect 1517 2904 1529 2944
rect 1537 2904 1549 2944
rect 1577 2904 1589 2944
rect 1599 2904 1611 2984
rect 1619 2904 1631 2984
rect 1662 2904 1674 2984
rect 1690 2904 1702 2984
rect 1712 2904 1724 2944
rect 1762 2904 1774 2984
rect 1790 2904 1802 2984
rect 1812 2904 1824 2944
rect 1857 2904 1869 2984
rect 1885 2904 1897 2984
rect 1937 2904 1949 2976
rect 1957 2904 1969 2972
rect 1977 2904 1989 2984
rect 1997 2904 2009 2984
rect 2037 2904 2049 2944
rect 2057 2904 2069 2944
rect 2102 2904 2114 2984
rect 2130 2904 2142 2984
rect 2152 2904 2164 2944
rect 2197 2904 2209 2984
rect 2225 2904 2237 2984
rect 2291 2904 2303 2944
rect 2311 2904 2323 2944
rect 2331 2904 2343 2944
rect 2362 2904 2374 2984
rect 2390 2904 2402 2984
rect 2412 2904 2424 2944
rect 2457 2904 2469 2944
rect 2477 2904 2489 2944
rect 2522 2904 2534 2984
rect 2550 2904 2562 2984
rect 2572 2904 2584 2944
rect 2617 2904 2629 2944
rect 2639 2904 2651 2984
rect 2659 2904 2671 2984
rect 2697 2904 2709 2944
rect 2717 2904 2729 2944
rect 2737 2904 2749 2944
rect 2781 2904 2793 2984
rect 2801 2904 2813 2944
rect 2835 2904 2847 2944
rect 2867 2904 2879 2944
rect 2887 2904 2899 2944
rect 2913 2904 2925 2944
rect 2941 2904 2953 2924
rect 2971 2904 2983 2924
rect 2991 2904 3003 2984
rect 3043 2904 3055 2984
rect 3071 2904 3083 2984
rect 3111 2904 3123 2984
rect 3131 2904 3143 2984
rect 3151 2904 3163 2972
rect 3171 2904 3183 2976
rect 3197 2904 3209 2984
rect 3225 2904 3237 2984
rect 3281 2904 3293 2984
rect 3301 2904 3313 2944
rect 3335 2904 3347 2944
rect 3367 2904 3379 2944
rect 3387 2904 3399 2944
rect 3413 2904 3425 2944
rect 3441 2904 3453 2924
rect 3471 2904 3483 2924
rect 3491 2904 3503 2984
rect 3521 2904 3533 2984
rect 3541 2904 3553 2944
rect 3575 2904 3587 2944
rect 3607 2904 3619 2944
rect 3627 2904 3639 2944
rect 3653 2904 3665 2944
rect 3681 2904 3693 2924
rect 3711 2904 3723 2924
rect 3731 2904 3743 2984
rect 3757 2904 3769 2984
rect 3785 2904 3797 2984
rect 3856 2904 3868 2944
rect 3878 2904 3890 2984
rect 3906 2904 3918 2984
rect 3956 2904 3968 2944
rect 3978 2904 3990 2984
rect 4006 2904 4018 2984
rect 4042 2904 4054 2984
rect 4070 2904 4082 2984
rect 4092 2904 4104 2944
rect 4142 2904 4154 2984
rect 4170 2904 4182 2984
rect 4192 2904 4204 2944
rect 4237 2904 4249 2944
rect 4257 2904 4269 2944
rect 4297 2904 4309 2944
rect 4317 2904 4329 2944
rect 4337 2904 4349 2940
rect 4357 2904 4369 2944
rect 4397 2904 4409 2984
rect 4417 2904 4429 2924
rect 4447 2904 4459 2924
rect 4475 2904 4487 2944
rect 4501 2904 4513 2944
rect 4521 2904 4533 2944
rect 4553 2904 4565 2944
rect 4587 2904 4599 2944
rect 4607 2904 4619 2984
rect 4642 2904 4654 2984
rect 4670 2904 4682 2984
rect 4692 2904 4704 2944
rect 31 2836 43 2876
rect 51 2836 63 2876
rect 96 2836 108 2876
rect 118 2796 130 2876
rect 146 2796 158 2876
rect 177 2798 189 2876
rect 197 2810 209 2876
rect 217 2798 229 2876
rect 237 2796 249 2864
rect 257 2796 269 2876
rect 297 2836 309 2876
rect 317 2836 329 2876
rect 337 2836 349 2876
rect 377 2836 389 2876
rect 397 2836 409 2876
rect 421 2796 433 2876
rect 441 2796 453 2876
rect 496 2836 508 2876
rect 518 2796 530 2876
rect 546 2796 558 2876
rect 577 2836 589 2876
rect 597 2836 609 2876
rect 617 2836 629 2876
rect 671 2796 683 2876
rect 691 2796 703 2876
rect 731 2796 743 2876
rect 751 2796 763 2876
rect 777 2836 789 2876
rect 797 2836 809 2876
rect 817 2836 829 2876
rect 857 2836 869 2876
rect 877 2836 889 2876
rect 901 2796 913 2876
rect 921 2796 933 2876
rect 976 2836 988 2876
rect 998 2796 1010 2876
rect 1026 2796 1038 2876
rect 1057 2836 1069 2876
rect 1077 2836 1089 2876
rect 1097 2836 1109 2876
rect 1156 2836 1168 2876
rect 1178 2796 1190 2876
rect 1206 2796 1218 2876
rect 1237 2796 1249 2876
rect 1257 2856 1269 2876
rect 1287 2856 1299 2876
rect 1315 2836 1327 2876
rect 1341 2836 1353 2876
rect 1361 2836 1373 2876
rect 1393 2836 1405 2876
rect 1427 2836 1439 2876
rect 1447 2796 1459 2876
rect 1489 2796 1501 2876
rect 1509 2796 1521 2876
rect 1531 2836 1543 2876
rect 1561 2796 1573 2876
rect 1581 2836 1593 2876
rect 1615 2836 1627 2876
rect 1647 2836 1659 2876
rect 1667 2836 1679 2876
rect 1693 2836 1705 2876
rect 1721 2856 1733 2876
rect 1751 2856 1763 2876
rect 1771 2796 1783 2876
rect 1802 2796 1814 2876
rect 1830 2796 1842 2876
rect 1852 2836 1864 2876
rect 1897 2836 1909 2876
rect 1917 2836 1929 2876
rect 1957 2796 1969 2876
rect 1987 2796 2009 2876
rect 2027 2796 2039 2876
rect 2103 2796 2115 2876
rect 2131 2796 2143 2876
rect 2183 2796 2195 2876
rect 2211 2796 2223 2876
rect 2263 2796 2275 2876
rect 2291 2796 2303 2876
rect 2317 2836 2329 2876
rect 2337 2836 2349 2876
rect 2403 2796 2415 2876
rect 2431 2796 2443 2876
rect 2457 2836 2469 2876
rect 2477 2836 2489 2876
rect 2517 2836 2529 2876
rect 2537 2836 2549 2876
rect 2561 2796 2573 2876
rect 2581 2796 2593 2876
rect 2622 2796 2634 2876
rect 2650 2796 2662 2876
rect 2672 2836 2684 2876
rect 2722 2796 2734 2876
rect 2750 2796 2762 2876
rect 2772 2836 2784 2876
rect 2817 2836 2829 2876
rect 2837 2836 2849 2876
rect 2857 2836 2869 2876
rect 2901 2796 2913 2876
rect 2921 2836 2933 2876
rect 2955 2836 2967 2876
rect 2987 2836 2999 2876
rect 3007 2836 3019 2876
rect 3033 2836 3045 2876
rect 3061 2856 3073 2876
rect 3091 2856 3103 2876
rect 3111 2796 3123 2876
rect 3141 2796 3153 2876
rect 3161 2836 3173 2876
rect 3195 2836 3207 2876
rect 3227 2836 3239 2876
rect 3247 2836 3259 2876
rect 3273 2836 3285 2876
rect 3301 2856 3313 2876
rect 3331 2856 3343 2876
rect 3351 2796 3363 2876
rect 3391 2836 3403 2876
rect 3411 2836 3423 2876
rect 3463 2796 3475 2876
rect 3491 2796 3503 2876
rect 3531 2796 3543 2876
rect 3551 2796 3563 2876
rect 3581 2796 3593 2876
rect 3601 2836 3613 2876
rect 3635 2836 3647 2876
rect 3667 2836 3679 2876
rect 3687 2836 3699 2876
rect 3713 2836 3725 2876
rect 3741 2856 3753 2876
rect 3771 2856 3783 2876
rect 3791 2796 3803 2876
rect 3831 2796 3843 2876
rect 3851 2796 3863 2864
rect 3871 2798 3883 2876
rect 3891 2810 3903 2876
rect 3911 2798 3923 2876
rect 3963 2796 3975 2876
rect 3991 2796 4003 2876
rect 4022 2796 4034 2876
rect 4050 2796 4062 2876
rect 4072 2836 4084 2876
rect 4136 2836 4148 2876
rect 4158 2796 4170 2876
rect 4186 2796 4198 2876
rect 4217 2796 4229 2876
rect 4245 2796 4257 2876
rect 4301 2796 4313 2876
rect 4321 2836 4333 2876
rect 4355 2836 4367 2876
rect 4387 2836 4399 2876
rect 4407 2836 4419 2876
rect 4433 2836 4445 2876
rect 4461 2856 4473 2876
rect 4491 2856 4503 2876
rect 4511 2796 4523 2876
rect 4542 2796 4554 2876
rect 4570 2796 4582 2876
rect 4592 2836 4604 2876
rect 4637 2836 4649 2876
rect 4657 2836 4669 2876
rect 4677 2836 4689 2876
rect 17 2424 29 2464
rect 37 2424 49 2464
rect 57 2424 69 2460
rect 77 2424 89 2464
rect 117 2424 129 2496
rect 137 2424 149 2492
rect 157 2424 169 2504
rect 177 2424 189 2504
rect 231 2424 243 2464
rect 251 2424 263 2464
rect 287 2424 299 2504
rect 307 2424 319 2504
rect 331 2424 343 2464
rect 351 2424 363 2464
rect 391 2424 403 2504
rect 411 2424 423 2504
rect 431 2424 443 2492
rect 451 2424 463 2496
rect 491 2424 503 2464
rect 511 2424 523 2460
rect 531 2424 543 2464
rect 551 2424 563 2464
rect 596 2424 608 2464
rect 618 2424 630 2504
rect 646 2424 658 2504
rect 691 2424 703 2504
rect 711 2424 723 2504
rect 751 2424 763 2464
rect 771 2424 783 2464
rect 791 2424 803 2464
rect 831 2424 843 2464
rect 851 2424 863 2460
rect 871 2424 883 2464
rect 891 2424 903 2464
rect 936 2424 948 2464
rect 958 2424 970 2504
rect 986 2424 998 2504
rect 1017 2424 1029 2464
rect 1037 2424 1049 2464
rect 1057 2424 1069 2464
rect 1111 2424 1123 2464
rect 1131 2424 1143 2460
rect 1151 2424 1163 2464
rect 1171 2424 1183 2464
rect 1211 2424 1223 2464
rect 1231 2424 1243 2464
rect 1276 2424 1288 2464
rect 1298 2424 1310 2504
rect 1326 2424 1338 2504
rect 1357 2424 1369 2464
rect 1377 2424 1389 2464
rect 1397 2424 1409 2464
rect 1437 2424 1449 2504
rect 1457 2424 1469 2504
rect 1511 2424 1523 2464
rect 1531 2424 1543 2464
rect 1551 2424 1563 2464
rect 1581 2424 1593 2504
rect 1601 2424 1613 2464
rect 1635 2424 1647 2464
rect 1667 2424 1679 2464
rect 1687 2424 1699 2464
rect 1713 2424 1725 2464
rect 1741 2424 1753 2444
rect 1771 2424 1783 2444
rect 1791 2424 1803 2504
rect 1817 2424 1829 2464
rect 1837 2424 1849 2464
rect 1857 2424 1869 2464
rect 1897 2424 1909 2464
rect 1917 2424 1929 2464
rect 1937 2424 1949 2464
rect 1977 2424 1989 2464
rect 1997 2424 2009 2464
rect 2017 2424 2029 2460
rect 2037 2424 2049 2464
rect 2077 2424 2089 2504
rect 2105 2424 2117 2504
rect 2171 2424 2183 2464
rect 2191 2424 2203 2464
rect 2243 2424 2255 2504
rect 2271 2424 2283 2504
rect 2311 2424 2323 2464
rect 2331 2424 2343 2464
rect 2376 2424 2388 2464
rect 2398 2424 2410 2504
rect 2426 2424 2438 2504
rect 2457 2424 2469 2504
rect 2485 2424 2497 2504
rect 2537 2424 2549 2464
rect 2557 2424 2569 2464
rect 2581 2424 2593 2504
rect 2601 2424 2613 2504
rect 2642 2424 2654 2504
rect 2670 2424 2682 2504
rect 2692 2424 2704 2464
rect 2751 2424 2763 2464
rect 2771 2424 2783 2464
rect 2791 2424 2803 2464
rect 2817 2424 2829 2504
rect 2847 2424 2859 2503
rect 2867 2424 2879 2503
rect 2917 2424 2929 2464
rect 2937 2424 2949 2464
rect 2957 2424 2969 2464
rect 2997 2424 3009 2464
rect 3019 2424 3031 2504
rect 3039 2424 3051 2504
rect 3082 2424 3094 2504
rect 3110 2424 3122 2504
rect 3132 2424 3144 2464
rect 3189 2424 3201 2504
rect 3209 2424 3221 2504
rect 3231 2424 3243 2464
rect 3271 2424 3283 2464
rect 3291 2424 3303 2464
rect 3311 2424 3323 2464
rect 3337 2424 3349 2502
rect 3357 2424 3369 2490
rect 3377 2424 3389 2502
rect 3397 2436 3409 2504
rect 3417 2424 3429 2504
rect 3457 2424 3469 2464
rect 3479 2424 3491 2504
rect 3499 2424 3511 2504
rect 3549 2424 3561 2504
rect 3569 2424 3581 2504
rect 3591 2424 3603 2464
rect 3621 2424 3633 2504
rect 3641 2424 3653 2464
rect 3675 2424 3687 2464
rect 3707 2424 3719 2464
rect 3727 2424 3739 2464
rect 3753 2424 3765 2464
rect 3781 2424 3793 2444
rect 3811 2424 3823 2444
rect 3831 2424 3843 2504
rect 3871 2424 3883 2504
rect 3891 2424 3903 2504
rect 3911 2424 3923 2492
rect 3931 2424 3943 2496
rect 3957 2424 3969 2504
rect 3985 2424 3997 2504
rect 4037 2424 4049 2504
rect 4057 2424 4069 2504
rect 4077 2424 4089 2504
rect 4097 2424 4109 2504
rect 4117 2424 4129 2504
rect 4137 2424 4149 2504
rect 4157 2424 4169 2504
rect 4177 2424 4189 2504
rect 4197 2424 4209 2504
rect 4241 2424 4253 2504
rect 4261 2424 4273 2464
rect 4295 2424 4307 2464
rect 4327 2424 4339 2464
rect 4347 2424 4359 2464
rect 4373 2424 4385 2464
rect 4401 2424 4413 2444
rect 4431 2424 4443 2444
rect 4451 2424 4463 2504
rect 4482 2424 4494 2504
rect 4510 2424 4522 2504
rect 4532 2424 4544 2464
rect 4577 2424 4589 2464
rect 4597 2424 4609 2464
rect 4617 2424 4629 2464
rect 4657 2424 4669 2464
rect 4677 2424 4689 2464
rect 4697 2424 4709 2464
rect 31 2356 43 2396
rect 51 2360 63 2396
rect 71 2356 83 2396
rect 91 2356 103 2396
rect 136 2356 148 2396
rect 158 2316 170 2396
rect 186 2316 198 2396
rect 222 2316 234 2396
rect 250 2316 262 2396
rect 272 2356 284 2396
rect 317 2356 329 2396
rect 337 2356 349 2396
rect 357 2360 369 2396
rect 377 2356 389 2396
rect 417 2324 429 2396
rect 437 2328 449 2396
rect 457 2316 469 2396
rect 477 2316 489 2396
rect 522 2316 534 2396
rect 550 2316 562 2396
rect 572 2356 584 2396
rect 631 2316 643 2396
rect 651 2316 663 2396
rect 671 2328 683 2396
rect 691 2324 703 2396
rect 717 2356 729 2396
rect 737 2356 749 2396
rect 787 2316 799 2396
rect 807 2316 819 2396
rect 831 2356 843 2396
rect 851 2356 863 2396
rect 877 2356 889 2396
rect 897 2356 909 2396
rect 917 2356 929 2396
rect 957 2356 969 2396
rect 977 2356 989 2396
rect 1001 2316 1013 2396
rect 1021 2316 1033 2396
rect 1076 2356 1088 2396
rect 1098 2316 1110 2396
rect 1126 2316 1138 2396
rect 1176 2356 1188 2396
rect 1198 2316 1210 2396
rect 1226 2316 1238 2396
rect 1261 2316 1273 2396
rect 1281 2356 1293 2396
rect 1315 2356 1327 2396
rect 1347 2356 1359 2396
rect 1367 2356 1379 2396
rect 1393 2356 1405 2396
rect 1421 2376 1433 2396
rect 1451 2376 1463 2396
rect 1471 2316 1483 2396
rect 1516 2356 1528 2396
rect 1538 2316 1550 2396
rect 1566 2316 1578 2396
rect 1601 2316 1613 2396
rect 1621 2356 1633 2396
rect 1655 2356 1667 2396
rect 1687 2356 1699 2396
rect 1707 2356 1719 2396
rect 1733 2356 1745 2396
rect 1761 2376 1773 2396
rect 1791 2376 1803 2396
rect 1811 2316 1823 2396
rect 1851 2356 1863 2396
rect 1871 2356 1883 2396
rect 1911 2356 1923 2396
rect 1931 2356 1943 2396
rect 1962 2316 1974 2396
rect 1990 2316 2002 2396
rect 2012 2356 2024 2396
rect 2061 2316 2073 2396
rect 2081 2356 2093 2396
rect 2115 2356 2127 2396
rect 2147 2356 2159 2396
rect 2167 2356 2179 2396
rect 2193 2356 2205 2396
rect 2221 2376 2233 2396
rect 2251 2376 2263 2396
rect 2271 2316 2283 2396
rect 2311 2316 2323 2396
rect 2331 2316 2343 2396
rect 2351 2328 2363 2396
rect 2371 2324 2383 2396
rect 2411 2316 2423 2396
rect 2431 2316 2443 2396
rect 2451 2328 2463 2396
rect 2471 2324 2483 2396
rect 2497 2356 2509 2396
rect 2517 2356 2529 2396
rect 2537 2360 2549 2396
rect 2557 2356 2569 2396
rect 2597 2356 2609 2396
rect 2617 2356 2629 2396
rect 2641 2316 2653 2396
rect 2661 2316 2673 2396
rect 2697 2316 2709 2396
rect 2717 2376 2729 2396
rect 2747 2376 2759 2396
rect 2775 2356 2787 2396
rect 2801 2356 2813 2396
rect 2821 2356 2833 2396
rect 2853 2356 2865 2396
rect 2887 2356 2899 2396
rect 2907 2316 2919 2396
rect 2956 2356 2968 2396
rect 2978 2316 2990 2396
rect 3006 2316 3018 2396
rect 3056 2356 3068 2396
rect 3078 2316 3090 2396
rect 3106 2316 3118 2396
rect 3142 2316 3154 2396
rect 3170 2316 3182 2396
rect 3192 2356 3204 2396
rect 3237 2316 3249 2396
rect 3257 2376 3269 2396
rect 3287 2376 3299 2396
rect 3315 2356 3327 2396
rect 3341 2356 3353 2396
rect 3361 2356 3373 2396
rect 3393 2356 3405 2396
rect 3427 2356 3439 2396
rect 3447 2316 3459 2396
rect 3496 2356 3508 2396
rect 3518 2316 3530 2396
rect 3546 2316 3558 2396
rect 3603 2316 3615 2396
rect 3631 2316 3643 2396
rect 3657 2316 3669 2396
rect 3687 2317 3699 2396
rect 3707 2317 3719 2396
rect 3771 2356 3783 2396
rect 3791 2356 3803 2396
rect 3811 2356 3823 2396
rect 3851 2316 3863 2396
rect 3871 2316 3883 2384
rect 3891 2318 3903 2396
rect 3911 2330 3923 2396
rect 3931 2318 3943 2396
rect 3971 2316 3983 2396
rect 3991 2316 4003 2384
rect 4011 2318 4023 2396
rect 4031 2330 4043 2396
rect 4051 2318 4063 2396
rect 4081 2316 4093 2396
rect 4101 2356 4113 2396
rect 4135 2356 4147 2396
rect 4167 2356 4179 2396
rect 4187 2356 4199 2396
rect 4213 2356 4225 2396
rect 4241 2376 4253 2396
rect 4271 2376 4283 2396
rect 4291 2316 4303 2396
rect 4317 2316 4329 2396
rect 4337 2376 4349 2396
rect 4367 2376 4379 2396
rect 4395 2356 4407 2396
rect 4421 2356 4433 2396
rect 4441 2356 4453 2396
rect 4473 2356 4485 2396
rect 4507 2356 4519 2396
rect 4527 2316 4539 2396
rect 4562 2316 4574 2396
rect 4590 2316 4602 2396
rect 4612 2356 4624 2396
rect 4657 2356 4669 2396
rect 4677 2356 4689 2396
rect 4697 2356 4709 2396
rect 29 1944 41 2024
rect 49 1944 61 2024
rect 71 1944 83 1984
rect 116 1944 128 1984
rect 138 1944 150 2024
rect 166 1944 178 2024
rect 211 1944 223 1984
rect 231 1944 243 1980
rect 251 1944 263 1984
rect 271 1944 283 1984
rect 297 1944 309 2016
rect 317 1944 329 2012
rect 337 1944 349 2024
rect 357 1944 369 2024
rect 397 1944 409 2016
rect 417 1944 429 2012
rect 437 1944 449 2024
rect 457 1944 469 2024
rect 497 1944 509 1984
rect 517 1944 529 1984
rect 537 1944 549 1980
rect 557 1944 569 1984
rect 597 1944 609 1984
rect 617 1944 629 1984
rect 637 1944 649 1980
rect 657 1944 669 1984
rect 697 1944 709 2016
rect 717 1944 729 2012
rect 737 1944 749 2024
rect 757 1944 769 2024
rect 816 1944 828 1984
rect 838 1944 850 2024
rect 866 1944 878 2024
rect 897 1944 909 1984
rect 917 1944 929 1984
rect 937 1944 949 1980
rect 957 1944 969 1984
rect 997 1944 1009 1984
rect 1017 1944 1029 1984
rect 1037 1944 1049 1980
rect 1057 1944 1069 1984
rect 1097 1944 1109 1984
rect 1117 1944 1129 1984
rect 1137 1944 1149 1980
rect 1157 1944 1169 1984
rect 1197 1944 1209 2016
rect 1217 1944 1229 2012
rect 1237 1944 1249 2024
rect 1257 1944 1269 2024
rect 1297 1944 1309 2024
rect 1325 1944 1337 2024
rect 1391 1944 1403 1984
rect 1411 1944 1423 1984
rect 1431 1944 1443 1984
rect 1471 1944 1483 1984
rect 1491 1944 1503 1984
rect 1511 1944 1523 1984
rect 1537 1944 1549 1984
rect 1557 1944 1569 1984
rect 1577 1944 1589 1984
rect 1636 1944 1648 1984
rect 1658 1944 1670 2024
rect 1686 1944 1698 2024
rect 1717 1944 1729 2016
rect 1737 1944 1749 2012
rect 1757 1944 1769 2024
rect 1777 1944 1789 2024
rect 1817 1944 1829 2024
rect 1845 1944 1857 2024
rect 1916 1944 1928 1984
rect 1938 1944 1950 2024
rect 1966 1944 1978 2024
rect 2002 1944 2014 2024
rect 2030 1944 2042 2024
rect 2052 1944 2064 1984
rect 2116 1944 2128 1984
rect 2138 1944 2150 2024
rect 2166 1944 2178 2024
rect 2211 1944 2223 2024
rect 2231 1944 2243 2024
rect 2251 1944 2263 2024
rect 2271 1944 2283 2024
rect 2291 1944 2303 2024
rect 2311 1944 2323 2024
rect 2331 1944 2343 2024
rect 2351 1944 2363 2024
rect 2371 1944 2383 2024
rect 2397 1944 2409 1984
rect 2417 1944 2429 1984
rect 2437 1944 2449 1984
rect 2487 1944 2499 2024
rect 2507 1944 2519 2024
rect 2531 1944 2543 1984
rect 2551 1944 2563 1984
rect 2577 1944 2589 2024
rect 2607 1944 2619 2023
rect 2627 1944 2639 2023
rect 2691 1944 2703 1984
rect 2711 1944 2723 1984
rect 2731 1944 2743 1984
rect 2757 1944 2769 1984
rect 2777 1944 2789 1984
rect 2797 1944 2809 1984
rect 2841 1944 2853 2024
rect 2861 1944 2873 1984
rect 2895 1944 2907 1984
rect 2927 1944 2939 1984
rect 2947 1944 2959 1984
rect 2973 1944 2985 1984
rect 3001 1944 3013 1964
rect 3031 1944 3043 1964
rect 3051 1944 3063 2024
rect 3091 1944 3103 2024
rect 3111 1944 3123 2024
rect 3131 1944 3143 2012
rect 3151 1944 3163 2016
rect 3177 1944 3189 2024
rect 3205 1944 3217 2024
rect 3271 1944 3283 2024
rect 3291 1956 3303 2024
rect 3311 1944 3323 2022
rect 3331 1944 3343 2010
rect 3351 1944 3363 2022
rect 3381 1944 3393 2024
rect 3401 1944 3413 1984
rect 3435 1944 3447 1984
rect 3467 1944 3479 1984
rect 3487 1944 3499 1984
rect 3513 1944 3525 1984
rect 3541 1944 3553 1964
rect 3571 1944 3583 1964
rect 3591 1944 3603 2024
rect 3622 1944 3634 2024
rect 3650 1944 3662 2024
rect 3672 1944 3684 1984
rect 3721 1944 3733 2024
rect 3741 1944 3753 1984
rect 3775 1944 3787 1984
rect 3807 1944 3819 1984
rect 3827 1944 3839 1984
rect 3853 1944 3865 1984
rect 3881 1944 3893 1964
rect 3911 1944 3923 1964
rect 3931 1944 3943 2024
rect 3957 1944 3969 2024
rect 3977 1944 3989 1964
rect 4007 1944 4019 1964
rect 4035 1944 4047 1984
rect 4061 1944 4073 1984
rect 4081 1944 4093 1984
rect 4113 1944 4125 1984
rect 4147 1944 4159 1984
rect 4167 1944 4179 2024
rect 4211 1944 4223 2024
rect 4231 1956 4243 2024
rect 4251 1944 4263 2022
rect 4271 1944 4283 2010
rect 4291 1944 4303 2022
rect 4317 1944 4329 1984
rect 4337 1944 4349 1984
rect 4403 1944 4415 2024
rect 4431 1944 4443 2024
rect 4483 1944 4495 2024
rect 4511 1944 4523 2024
rect 4537 1944 4549 2024
rect 4557 1944 4569 1964
rect 4587 1944 4599 1964
rect 4615 1944 4627 1984
rect 4641 1944 4653 1984
rect 4661 1944 4673 1984
rect 4693 1944 4705 1984
rect 4727 1944 4739 1984
rect 4747 1944 4759 2024
rect 31 1836 43 1916
rect 51 1836 63 1904
rect 71 1838 83 1916
rect 91 1850 103 1916
rect 111 1838 123 1916
rect 142 1836 154 1916
rect 170 1836 182 1916
rect 192 1876 204 1916
rect 237 1876 249 1916
rect 257 1876 269 1916
rect 277 1876 289 1916
rect 331 1876 343 1916
rect 351 1880 363 1916
rect 371 1876 383 1916
rect 391 1876 403 1916
rect 417 1838 429 1916
rect 437 1850 449 1916
rect 457 1838 469 1916
rect 477 1836 489 1904
rect 497 1836 509 1916
rect 537 1876 549 1916
rect 557 1876 569 1916
rect 581 1836 593 1916
rect 601 1836 613 1916
rect 651 1836 663 1916
rect 671 1836 683 1916
rect 697 1876 709 1916
rect 719 1836 731 1916
rect 739 1836 751 1916
rect 796 1876 808 1916
rect 818 1836 830 1916
rect 846 1836 858 1916
rect 882 1836 894 1916
rect 910 1836 922 1916
rect 932 1876 944 1916
rect 977 1876 989 1916
rect 997 1876 1009 1916
rect 1017 1880 1029 1916
rect 1037 1876 1049 1916
rect 1077 1876 1089 1916
rect 1097 1876 1109 1916
rect 1137 1876 1149 1916
rect 1157 1876 1169 1916
rect 1177 1880 1189 1916
rect 1197 1876 1209 1916
rect 1237 1876 1249 1916
rect 1257 1876 1269 1916
rect 1277 1880 1289 1916
rect 1297 1876 1309 1916
rect 1351 1876 1363 1916
rect 1371 1876 1383 1916
rect 1411 1836 1423 1916
rect 1431 1836 1443 1904
rect 1451 1838 1463 1916
rect 1471 1850 1483 1916
rect 1491 1838 1503 1916
rect 1517 1876 1529 1916
rect 1537 1876 1549 1916
rect 1557 1880 1569 1916
rect 1577 1876 1589 1916
rect 1617 1876 1629 1916
rect 1637 1876 1649 1916
rect 1691 1836 1703 1916
rect 1711 1836 1723 1916
rect 1751 1876 1763 1916
rect 1771 1880 1783 1916
rect 1791 1876 1803 1916
rect 1811 1876 1823 1916
rect 1837 1876 1849 1916
rect 1857 1876 1869 1916
rect 1881 1836 1893 1916
rect 1901 1836 1913 1916
rect 1941 1836 1953 1916
rect 1961 1876 1973 1916
rect 1995 1876 2007 1916
rect 2027 1876 2039 1916
rect 2047 1876 2059 1916
rect 2073 1876 2085 1916
rect 2101 1896 2113 1916
rect 2131 1896 2143 1916
rect 2151 1836 2163 1916
rect 2203 1836 2215 1916
rect 2231 1836 2243 1916
rect 2257 1876 2269 1916
rect 2277 1876 2289 1916
rect 2322 1836 2334 1916
rect 2350 1836 2362 1916
rect 2372 1876 2384 1916
rect 2417 1836 2429 1916
rect 2445 1836 2457 1916
rect 2497 1836 2509 1916
rect 2525 1836 2537 1916
rect 2582 1836 2594 1916
rect 2610 1836 2622 1916
rect 2632 1876 2644 1916
rect 2691 1876 2703 1916
rect 2711 1876 2723 1916
rect 2731 1876 2743 1916
rect 2783 1836 2795 1916
rect 2811 1836 2823 1916
rect 2842 1836 2854 1916
rect 2870 1836 2882 1916
rect 2892 1876 2904 1916
rect 2937 1876 2949 1916
rect 2957 1876 2969 1916
rect 3023 1836 3035 1916
rect 3051 1836 3063 1916
rect 3077 1836 3089 1916
rect 3097 1896 3109 1916
rect 3127 1896 3139 1916
rect 3155 1876 3167 1916
rect 3181 1876 3193 1916
rect 3201 1876 3213 1916
rect 3233 1876 3245 1916
rect 3267 1876 3279 1916
rect 3287 1836 3299 1916
rect 3322 1836 3334 1916
rect 3350 1836 3362 1916
rect 3372 1876 3384 1916
rect 3417 1876 3429 1916
rect 3437 1876 3449 1916
rect 3457 1876 3469 1916
rect 3497 1836 3509 1916
rect 3517 1896 3529 1916
rect 3547 1896 3559 1916
rect 3575 1876 3587 1916
rect 3601 1876 3613 1916
rect 3621 1876 3633 1916
rect 3653 1876 3665 1916
rect 3687 1876 3699 1916
rect 3707 1836 3719 1916
rect 3737 1876 3749 1916
rect 3759 1836 3771 1916
rect 3779 1836 3791 1916
rect 3831 1876 3843 1916
rect 3851 1876 3863 1916
rect 3871 1876 3883 1916
rect 3916 1876 3928 1916
rect 3938 1836 3950 1916
rect 3966 1836 3978 1916
rect 4016 1876 4028 1916
rect 4038 1836 4050 1916
rect 4066 1836 4078 1916
rect 4097 1836 4109 1916
rect 4127 1837 4139 1916
rect 4147 1837 4159 1916
rect 4211 1876 4223 1916
rect 4231 1876 4243 1916
rect 4257 1844 4269 1916
rect 4277 1848 4289 1916
rect 4297 1836 4309 1916
rect 4317 1836 4329 1916
rect 4383 1836 4395 1916
rect 4411 1836 4423 1916
rect 4437 1836 4449 1916
rect 4457 1896 4469 1916
rect 4487 1896 4499 1916
rect 4515 1876 4527 1916
rect 4541 1876 4553 1916
rect 4561 1876 4573 1916
rect 4593 1876 4605 1916
rect 4627 1876 4639 1916
rect 4647 1836 4659 1916
rect 4691 1876 4703 1916
rect 4711 1876 4723 1916
rect 4731 1876 4743 1916
rect 31 1464 43 1504
rect 51 1464 63 1504
rect 91 1464 103 1544
rect 111 1464 123 1544
rect 131 1464 143 1532
rect 151 1464 163 1536
rect 177 1464 189 1504
rect 197 1464 209 1504
rect 217 1464 229 1500
rect 237 1464 249 1504
rect 277 1464 289 1504
rect 297 1464 309 1504
rect 317 1464 329 1504
rect 376 1464 388 1504
rect 398 1464 410 1544
rect 426 1464 438 1544
rect 469 1464 481 1544
rect 489 1464 501 1544
rect 511 1464 523 1504
rect 551 1464 563 1504
rect 571 1464 583 1504
rect 597 1464 609 1504
rect 617 1464 629 1504
rect 637 1464 649 1500
rect 657 1464 669 1504
rect 697 1464 709 1536
rect 717 1464 729 1532
rect 737 1464 749 1544
rect 757 1464 769 1544
rect 797 1464 809 1504
rect 817 1464 829 1504
rect 837 1464 849 1500
rect 857 1464 869 1504
rect 897 1464 909 1536
rect 917 1464 929 1532
rect 937 1464 949 1544
rect 957 1464 969 1544
rect 997 1464 1009 1504
rect 1017 1464 1029 1504
rect 1037 1464 1049 1500
rect 1057 1464 1069 1504
rect 1116 1464 1128 1504
rect 1138 1464 1150 1544
rect 1166 1464 1178 1544
rect 1197 1464 1209 1504
rect 1217 1464 1229 1504
rect 1237 1464 1249 1500
rect 1257 1464 1269 1504
rect 1297 1464 1309 1536
rect 1317 1464 1329 1532
rect 1337 1464 1349 1544
rect 1357 1464 1369 1544
rect 1411 1464 1423 1504
rect 1431 1464 1443 1504
rect 1457 1464 1469 1504
rect 1477 1464 1489 1504
rect 1497 1464 1509 1500
rect 1517 1464 1529 1504
rect 1557 1464 1569 1536
rect 1577 1464 1589 1532
rect 1597 1464 1609 1544
rect 1617 1464 1629 1544
rect 1657 1464 1669 1504
rect 1677 1464 1689 1504
rect 1697 1464 1709 1500
rect 1717 1464 1729 1504
rect 1762 1464 1774 1544
rect 1790 1464 1802 1544
rect 1812 1464 1824 1504
rect 1871 1464 1883 1544
rect 1891 1464 1903 1544
rect 1911 1464 1923 1532
rect 1931 1464 1943 1536
rect 1957 1464 1969 1504
rect 1977 1464 1989 1504
rect 2017 1464 2029 1504
rect 2037 1464 2049 1504
rect 2057 1464 2069 1500
rect 2077 1464 2089 1504
rect 2136 1464 2148 1504
rect 2158 1464 2170 1544
rect 2186 1464 2198 1544
rect 2217 1464 2229 1504
rect 2237 1464 2249 1504
rect 2277 1464 2289 1544
rect 2297 1464 2309 1484
rect 2327 1464 2339 1484
rect 2355 1464 2367 1504
rect 2381 1464 2393 1504
rect 2401 1464 2413 1504
rect 2433 1464 2445 1504
rect 2467 1464 2479 1504
rect 2487 1464 2499 1544
rect 2536 1464 2548 1504
rect 2558 1464 2570 1544
rect 2586 1464 2598 1544
rect 2627 1464 2639 1544
rect 2647 1464 2659 1544
rect 2671 1464 2683 1504
rect 2691 1464 2703 1504
rect 2717 1464 2729 1544
rect 2745 1464 2757 1544
rect 2797 1464 2809 1536
rect 2817 1464 2829 1532
rect 2837 1464 2849 1544
rect 2857 1464 2869 1544
rect 2923 1464 2935 1544
rect 2951 1464 2963 1544
rect 2991 1464 3003 1504
rect 3011 1464 3023 1504
rect 3051 1464 3063 1504
rect 3071 1464 3083 1504
rect 3102 1464 3114 1544
rect 3130 1464 3142 1544
rect 3152 1464 3164 1504
rect 3197 1464 3209 1504
rect 3217 1464 3229 1504
rect 3237 1464 3249 1504
rect 3291 1464 3303 1504
rect 3311 1464 3323 1504
rect 3331 1464 3343 1504
rect 3376 1464 3388 1504
rect 3398 1464 3410 1544
rect 3426 1464 3438 1544
rect 3461 1464 3473 1544
rect 3481 1464 3493 1504
rect 3515 1464 3527 1504
rect 3547 1464 3559 1504
rect 3567 1464 3579 1504
rect 3593 1464 3605 1504
rect 3621 1464 3633 1484
rect 3651 1464 3663 1484
rect 3671 1464 3683 1544
rect 3697 1464 3709 1504
rect 3717 1464 3729 1504
rect 3771 1464 3783 1504
rect 3791 1464 3803 1504
rect 3836 1464 3848 1504
rect 3858 1464 3870 1544
rect 3886 1464 3898 1544
rect 3917 1464 3929 1544
rect 3945 1464 3957 1544
rect 3997 1464 4009 1544
rect 4025 1464 4037 1544
rect 4077 1464 4089 1504
rect 4097 1464 4109 1504
rect 4137 1464 4149 1536
rect 4157 1464 4169 1532
rect 4177 1464 4189 1544
rect 4197 1464 4209 1544
rect 4237 1464 4249 1544
rect 4265 1464 4277 1544
rect 4317 1464 4329 1536
rect 4337 1464 4349 1532
rect 4357 1464 4369 1544
rect 4377 1464 4389 1544
rect 4417 1464 4429 1504
rect 4437 1464 4449 1504
rect 4477 1464 4489 1504
rect 4497 1464 4509 1504
rect 4551 1464 4563 1504
rect 4571 1464 4583 1504
rect 4602 1464 4614 1544
rect 4630 1464 4642 1544
rect 4652 1464 4664 1504
rect 4697 1464 4709 1504
rect 4717 1464 4729 1504
rect 4737 1464 4749 1504
rect 31 1356 43 1436
rect 51 1356 63 1436
rect 71 1368 83 1436
rect 91 1364 103 1436
rect 117 1396 129 1436
rect 137 1396 149 1436
rect 157 1400 169 1436
rect 177 1396 189 1436
rect 217 1396 229 1436
rect 237 1396 249 1436
rect 257 1400 269 1436
rect 277 1396 289 1436
rect 331 1396 343 1436
rect 351 1396 363 1436
rect 371 1396 383 1436
rect 402 1356 414 1436
rect 430 1356 442 1436
rect 452 1396 464 1436
rect 497 1364 509 1436
rect 517 1368 529 1436
rect 537 1356 549 1436
rect 557 1356 569 1436
rect 602 1356 614 1436
rect 630 1356 642 1436
rect 652 1396 664 1436
rect 702 1356 714 1436
rect 730 1356 742 1436
rect 752 1396 764 1436
rect 797 1396 809 1436
rect 817 1396 829 1436
rect 841 1356 853 1436
rect 861 1356 873 1436
rect 911 1396 923 1436
rect 931 1396 943 1436
rect 951 1396 963 1436
rect 977 1396 989 1436
rect 997 1396 1009 1436
rect 1017 1396 1029 1436
rect 1071 1396 1083 1436
rect 1091 1400 1103 1436
rect 1111 1396 1123 1436
rect 1131 1396 1143 1436
rect 1171 1396 1183 1436
rect 1191 1396 1203 1436
rect 1227 1356 1239 1436
rect 1247 1356 1259 1436
rect 1271 1396 1283 1436
rect 1291 1396 1303 1436
rect 1322 1356 1334 1436
rect 1350 1356 1362 1436
rect 1372 1396 1384 1436
rect 1436 1396 1448 1436
rect 1458 1356 1470 1436
rect 1486 1356 1498 1436
rect 1517 1396 1529 1436
rect 1537 1396 1549 1436
rect 1557 1396 1569 1436
rect 1602 1356 1614 1436
rect 1630 1356 1642 1436
rect 1652 1396 1664 1436
rect 1697 1396 1709 1436
rect 1717 1396 1729 1436
rect 1737 1396 1749 1436
rect 1777 1364 1789 1436
rect 1797 1368 1809 1436
rect 1817 1356 1829 1436
rect 1837 1356 1849 1436
rect 1877 1396 1889 1436
rect 1897 1396 1909 1436
rect 1917 1400 1929 1436
rect 1937 1396 1949 1436
rect 1982 1356 1994 1436
rect 2010 1356 2022 1436
rect 2032 1396 2044 1436
rect 2077 1396 2089 1436
rect 2097 1396 2109 1436
rect 2137 1396 2149 1436
rect 2157 1396 2169 1436
rect 2177 1400 2189 1436
rect 2197 1396 2209 1436
rect 2237 1396 2249 1436
rect 2257 1396 2269 1436
rect 2277 1396 2289 1436
rect 2317 1356 2329 1436
rect 2347 1357 2359 1436
rect 2367 1357 2379 1436
rect 2431 1396 2443 1436
rect 2451 1396 2463 1436
rect 2471 1396 2483 1436
rect 2497 1396 2509 1436
rect 2517 1396 2529 1436
rect 2569 1356 2581 1436
rect 2589 1356 2601 1436
rect 2611 1396 2623 1436
rect 2642 1356 2654 1436
rect 2670 1356 2682 1436
rect 2692 1396 2704 1436
rect 2761 1356 2773 1436
rect 2791 1356 2813 1436
rect 2831 1356 2843 1436
rect 2861 1356 2873 1436
rect 2881 1396 2893 1436
rect 2915 1396 2927 1436
rect 2947 1396 2959 1436
rect 2967 1396 2979 1436
rect 2993 1396 3005 1436
rect 3021 1416 3033 1436
rect 3051 1416 3063 1436
rect 3071 1356 3083 1436
rect 3123 1356 3135 1436
rect 3151 1356 3163 1436
rect 3191 1356 3203 1436
rect 3211 1356 3223 1436
rect 3231 1368 3243 1436
rect 3251 1364 3263 1436
rect 3281 1356 3293 1436
rect 3301 1396 3313 1436
rect 3335 1396 3347 1436
rect 3367 1396 3379 1436
rect 3387 1396 3399 1436
rect 3413 1396 3425 1436
rect 3441 1416 3453 1436
rect 3471 1416 3483 1436
rect 3491 1356 3503 1436
rect 3531 1396 3543 1436
rect 3551 1396 3563 1436
rect 3603 1356 3615 1436
rect 3631 1356 3643 1436
rect 3683 1356 3695 1436
rect 3711 1356 3723 1436
rect 3737 1396 3749 1436
rect 3757 1396 3769 1436
rect 3797 1356 3809 1436
rect 3817 1416 3829 1436
rect 3847 1416 3859 1436
rect 3875 1396 3887 1436
rect 3901 1396 3913 1436
rect 3921 1396 3933 1436
rect 3953 1396 3965 1436
rect 3987 1396 3999 1436
rect 4007 1356 4019 1436
rect 4042 1356 4054 1436
rect 4070 1356 4082 1436
rect 4092 1396 4104 1436
rect 4137 1396 4149 1436
rect 4157 1396 4169 1436
rect 4177 1396 4189 1436
rect 4229 1356 4241 1436
rect 4249 1356 4261 1436
rect 4271 1396 4283 1436
rect 4311 1396 4323 1436
rect 4331 1396 4343 1436
rect 4351 1396 4363 1436
rect 4396 1396 4408 1436
rect 4418 1356 4430 1436
rect 4446 1356 4458 1436
rect 4496 1396 4508 1436
rect 4518 1356 4530 1436
rect 4546 1356 4558 1436
rect 4577 1356 4589 1436
rect 4605 1356 4617 1436
rect 4657 1396 4669 1436
rect 4677 1396 4689 1436
rect 4731 1396 4743 1436
rect 4751 1396 4763 1436
rect 36 984 48 1024
rect 58 984 70 1064
rect 86 984 98 1064
rect 122 984 134 1064
rect 150 984 162 1064
rect 172 984 184 1024
rect 217 984 229 1024
rect 237 984 249 1024
rect 257 984 269 1020
rect 277 984 289 1024
rect 317 984 329 1056
rect 337 984 349 1052
rect 357 984 369 1064
rect 377 984 389 1064
rect 417 984 429 1024
rect 437 984 449 1024
rect 457 984 469 1020
rect 477 984 489 1024
rect 517 984 529 1056
rect 537 984 549 1052
rect 557 984 569 1064
rect 577 984 589 1064
rect 631 984 643 1024
rect 651 984 663 1024
rect 671 984 683 1024
rect 707 984 719 1064
rect 727 984 739 1064
rect 751 984 763 1024
rect 771 984 783 1024
rect 811 984 823 1024
rect 831 984 843 1020
rect 851 984 863 1024
rect 871 984 883 1024
rect 916 984 928 1024
rect 938 984 950 1064
rect 966 984 978 1064
rect 1002 984 1014 1064
rect 1030 984 1042 1064
rect 1052 984 1064 1024
rect 1116 984 1128 1024
rect 1138 984 1150 1064
rect 1166 984 1178 1064
rect 1211 984 1223 1024
rect 1231 984 1243 1024
rect 1251 984 1263 1024
rect 1287 984 1299 1064
rect 1307 984 1319 1064
rect 1331 984 1343 1024
rect 1351 984 1363 1024
rect 1377 984 1389 1024
rect 1397 984 1409 1024
rect 1417 984 1429 1024
rect 1471 984 1483 1064
rect 1491 984 1503 1064
rect 1531 984 1543 1024
rect 1551 984 1563 1024
rect 1571 984 1583 1024
rect 1611 984 1623 1024
rect 1631 984 1643 1024
rect 1651 984 1663 1024
rect 1677 984 1689 1024
rect 1697 984 1709 1024
rect 1717 984 1729 1020
rect 1737 984 1749 1024
rect 1791 984 1803 1024
rect 1811 984 1823 1024
rect 1831 984 1843 1024
rect 1857 984 1869 1024
rect 1877 984 1889 1024
rect 1897 984 1909 1020
rect 1917 984 1929 1024
rect 1957 984 1969 1024
rect 1977 984 1989 1024
rect 1997 984 2009 1024
rect 2051 984 2063 1064
rect 2071 996 2083 1064
rect 2091 984 2103 1062
rect 2111 984 2123 1050
rect 2131 984 2143 1062
rect 2171 984 2183 1024
rect 2191 984 2203 1020
rect 2211 984 2223 1024
rect 2231 984 2243 1024
rect 2271 984 2283 1024
rect 2291 984 2303 1024
rect 2311 984 2323 1024
rect 2337 984 2349 1056
rect 2357 984 2369 1052
rect 2377 984 2389 1064
rect 2397 984 2409 1064
rect 2451 984 2463 1024
rect 2471 984 2483 1024
rect 2511 984 2523 1024
rect 2531 984 2543 1024
rect 2551 984 2563 1024
rect 2601 984 2613 1064
rect 2631 984 2653 1064
rect 2671 984 2683 1064
rect 2697 984 2709 1024
rect 2719 984 2731 1064
rect 2739 984 2751 1064
rect 2781 984 2793 1064
rect 2801 984 2813 1024
rect 2835 984 2847 1024
rect 2867 984 2879 1024
rect 2887 984 2899 1024
rect 2913 984 2925 1024
rect 2941 984 2953 1004
rect 2971 984 2983 1004
rect 2991 984 3003 1064
rect 3017 984 3029 1024
rect 3037 984 3049 1024
rect 3057 984 3069 1024
rect 3116 984 3128 1024
rect 3138 984 3150 1064
rect 3166 984 3178 1064
rect 3197 984 3209 1064
rect 3217 984 3229 1064
rect 3237 984 3249 1064
rect 3257 984 3269 1064
rect 3277 984 3289 1064
rect 3329 984 3341 1064
rect 3349 984 3361 1064
rect 3371 984 3383 1024
rect 3397 984 3409 1024
rect 3419 984 3431 1064
rect 3439 984 3451 1064
rect 3477 984 3489 1064
rect 3497 984 3509 1064
rect 3517 984 3529 1064
rect 3537 984 3549 1064
rect 3557 984 3569 1064
rect 3577 984 3589 1064
rect 3597 984 3609 1064
rect 3617 984 3629 1064
rect 3637 984 3649 1064
rect 3677 984 3689 1064
rect 3697 984 3709 1064
rect 3717 984 3729 1064
rect 3737 984 3749 1064
rect 3757 984 3769 1064
rect 3777 984 3789 1064
rect 3797 984 3809 1064
rect 3817 984 3829 1064
rect 3837 984 3849 1064
rect 3877 984 3889 1024
rect 3899 984 3911 1064
rect 3919 984 3931 1064
rect 3957 984 3969 1024
rect 3977 984 3989 1024
rect 3997 984 4009 1024
rect 4037 984 4049 1064
rect 4057 984 4069 1004
rect 4087 984 4099 1004
rect 4115 984 4127 1024
rect 4141 984 4153 1024
rect 4161 984 4173 1024
rect 4193 984 4205 1024
rect 4227 984 4239 1024
rect 4247 984 4259 1064
rect 4277 984 4289 1024
rect 4297 984 4309 1024
rect 4317 984 4329 1024
rect 4362 984 4374 1064
rect 4390 984 4402 1064
rect 4412 984 4424 1024
rect 4471 984 4483 1024
rect 4491 984 4503 1024
rect 4511 984 4523 1024
rect 4542 984 4554 1064
rect 4570 984 4582 1064
rect 4592 984 4604 1024
rect 4637 984 4649 1024
rect 4657 984 4669 1024
rect 4677 984 4689 1020
rect 4697 984 4709 1024
rect 31 916 43 956
rect 51 916 63 956
rect 71 916 83 956
rect 107 876 119 956
rect 127 876 139 956
rect 151 916 163 956
rect 171 916 183 956
rect 216 916 228 956
rect 238 876 250 956
rect 266 876 278 956
rect 311 876 323 956
rect 331 876 343 944
rect 351 878 363 956
rect 371 890 383 956
rect 391 878 403 956
rect 429 876 441 956
rect 449 876 461 956
rect 471 916 483 956
rect 497 916 509 956
rect 517 916 529 956
rect 571 916 583 956
rect 591 916 603 956
rect 631 876 643 956
rect 651 876 663 956
rect 671 888 683 956
rect 691 884 703 956
rect 717 916 729 956
rect 737 916 749 956
rect 757 920 769 956
rect 777 916 789 956
rect 827 876 839 956
rect 847 876 859 956
rect 871 916 883 956
rect 891 916 903 956
rect 917 916 929 956
rect 937 916 949 956
rect 957 916 969 956
rect 1011 916 1023 956
rect 1031 920 1043 956
rect 1051 916 1063 956
rect 1071 916 1083 956
rect 1102 876 1114 956
rect 1130 876 1142 956
rect 1152 916 1164 956
rect 1211 916 1223 956
rect 1231 920 1243 956
rect 1251 916 1263 956
rect 1271 916 1283 956
rect 1297 916 1309 956
rect 1317 916 1329 956
rect 1362 876 1374 956
rect 1390 876 1402 956
rect 1412 916 1424 956
rect 1471 916 1483 956
rect 1491 916 1503 956
rect 1511 916 1523 956
rect 1537 916 1549 956
rect 1557 916 1569 956
rect 1577 916 1589 956
rect 1636 916 1648 956
rect 1658 876 1670 956
rect 1686 876 1698 956
rect 1717 916 1729 956
rect 1737 916 1749 956
rect 1761 876 1773 956
rect 1781 876 1793 956
rect 1831 916 1843 956
rect 1851 916 1863 956
rect 1891 916 1903 956
rect 1911 916 1923 956
rect 1931 916 1943 956
rect 1957 916 1969 956
rect 1977 916 1989 956
rect 2031 916 2043 956
rect 2051 920 2063 956
rect 2071 916 2083 956
rect 2091 916 2103 956
rect 2117 916 2129 956
rect 2137 916 2149 956
rect 2182 876 2194 956
rect 2210 876 2222 956
rect 2232 916 2244 956
rect 2291 876 2303 956
rect 2311 876 2323 956
rect 2331 888 2343 956
rect 2351 884 2363 956
rect 2377 916 2389 956
rect 2397 916 2409 956
rect 2437 916 2449 956
rect 2457 916 2469 956
rect 2477 920 2489 956
rect 2497 916 2509 956
rect 2551 916 2563 956
rect 2571 920 2583 956
rect 2591 916 2603 956
rect 2611 916 2623 956
rect 2637 884 2649 956
rect 2657 888 2669 956
rect 2677 876 2689 956
rect 2697 876 2709 956
rect 2751 916 2763 956
rect 2771 916 2783 956
rect 2791 916 2803 956
rect 2841 876 2853 956
rect 2871 876 2893 956
rect 2911 876 2923 956
rect 2951 916 2963 956
rect 2971 916 2983 956
rect 3023 876 3035 956
rect 3051 876 3063 956
rect 3103 876 3115 956
rect 3131 876 3143 956
rect 3157 916 3169 956
rect 3177 916 3189 956
rect 3222 876 3234 956
rect 3250 876 3262 956
rect 3272 916 3284 956
rect 3317 916 3329 956
rect 3337 916 3349 956
rect 3357 916 3369 956
rect 3397 876 3409 956
rect 3417 936 3429 956
rect 3447 936 3459 956
rect 3475 916 3487 956
rect 3501 916 3513 956
rect 3521 916 3533 956
rect 3553 916 3565 956
rect 3587 916 3599 956
rect 3607 876 3619 956
rect 3637 916 3649 956
rect 3659 876 3671 956
rect 3679 876 3691 956
rect 3721 876 3733 956
rect 3741 916 3753 956
rect 3775 916 3787 956
rect 3807 916 3819 956
rect 3827 916 3839 956
rect 3853 916 3865 956
rect 3881 936 3893 956
rect 3911 936 3923 956
rect 3931 876 3943 956
rect 3976 916 3988 956
rect 3998 876 4010 956
rect 4026 876 4038 956
rect 4057 876 4069 956
rect 4077 936 4089 956
rect 4107 936 4119 956
rect 4135 916 4147 956
rect 4161 916 4173 956
rect 4181 916 4193 956
rect 4213 916 4225 956
rect 4247 916 4259 956
rect 4267 876 4279 956
rect 4301 876 4313 956
rect 4321 916 4333 956
rect 4355 916 4367 956
rect 4387 916 4399 956
rect 4407 916 4419 956
rect 4433 916 4445 956
rect 4461 936 4473 956
rect 4491 936 4503 956
rect 4511 876 4523 956
rect 4542 876 4554 956
rect 4570 876 4582 956
rect 4592 916 4604 956
rect 4642 876 4654 956
rect 4670 876 4682 956
rect 4692 916 4704 956
rect 43 504 55 584
rect 71 504 83 584
rect 111 504 123 584
rect 131 504 143 584
rect 151 504 163 572
rect 171 504 183 576
rect 197 504 209 544
rect 217 504 229 544
rect 271 504 283 584
rect 291 504 303 584
rect 311 504 323 572
rect 331 504 343 576
rect 357 504 369 544
rect 377 504 389 544
rect 397 504 409 540
rect 417 504 429 544
rect 476 504 488 544
rect 498 504 510 584
rect 526 504 538 584
rect 569 504 581 584
rect 589 504 601 584
rect 611 504 623 544
rect 656 504 668 544
rect 678 504 690 584
rect 706 504 718 584
rect 749 504 761 584
rect 769 504 781 584
rect 791 504 803 544
rect 817 504 829 544
rect 837 504 849 544
rect 861 504 873 584
rect 881 504 893 584
rect 922 504 934 584
rect 950 504 962 584
rect 972 504 984 544
rect 1036 504 1048 544
rect 1058 504 1070 584
rect 1086 504 1098 584
rect 1131 504 1143 584
rect 1151 504 1163 584
rect 1177 504 1189 576
rect 1197 504 1209 572
rect 1217 504 1229 584
rect 1237 504 1249 584
rect 1291 504 1303 544
rect 1311 504 1323 544
rect 1342 504 1354 584
rect 1370 504 1382 584
rect 1392 504 1404 544
rect 1442 504 1454 584
rect 1470 504 1482 584
rect 1492 504 1504 544
rect 1551 504 1563 584
rect 1571 504 1583 584
rect 1591 504 1603 572
rect 1611 504 1623 576
rect 1637 504 1649 576
rect 1657 504 1669 572
rect 1677 504 1689 584
rect 1697 504 1709 584
rect 1737 504 1749 544
rect 1757 504 1769 544
rect 1777 504 1789 540
rect 1797 504 1809 544
rect 1842 504 1854 584
rect 1870 504 1882 584
rect 1892 504 1904 544
rect 1951 504 1963 584
rect 1971 504 1983 584
rect 1991 504 2003 572
rect 2011 504 2023 576
rect 2042 504 2054 584
rect 2070 504 2082 584
rect 2092 504 2104 544
rect 2151 504 2163 544
rect 2171 504 2183 540
rect 2191 504 2203 544
rect 2211 504 2223 544
rect 2256 504 2268 544
rect 2278 504 2290 584
rect 2306 504 2318 584
rect 2342 504 2354 584
rect 2370 504 2382 584
rect 2392 504 2404 544
rect 2437 504 2449 544
rect 2457 504 2469 544
rect 2477 504 2489 540
rect 2497 504 2509 544
rect 2537 504 2549 544
rect 2557 504 2569 544
rect 2577 504 2589 540
rect 2597 504 2609 544
rect 2651 504 2663 544
rect 2671 504 2683 544
rect 2697 504 2709 544
rect 2717 504 2729 544
rect 2737 504 2749 540
rect 2757 504 2769 544
rect 2801 504 2813 584
rect 2821 504 2833 544
rect 2855 504 2867 544
rect 2887 504 2899 544
rect 2907 504 2919 544
rect 2933 504 2945 544
rect 2961 504 2973 524
rect 2991 504 3003 524
rect 3011 504 3023 584
rect 3042 504 3054 584
rect 3070 504 3082 584
rect 3092 504 3104 544
rect 3137 504 3149 544
rect 3157 504 3169 544
rect 3197 504 3209 544
rect 3217 504 3229 544
rect 3257 504 3269 544
rect 3277 504 3289 544
rect 3297 504 3309 540
rect 3317 504 3329 544
rect 3371 504 3383 544
rect 3391 504 3403 544
rect 3431 504 3443 544
rect 3451 504 3463 544
rect 3471 504 3483 544
rect 3516 504 3528 544
rect 3538 504 3550 584
rect 3566 504 3578 584
rect 3601 504 3613 584
rect 3621 504 3633 544
rect 3655 504 3667 544
rect 3687 504 3699 544
rect 3707 504 3719 544
rect 3733 504 3745 544
rect 3761 504 3773 524
rect 3791 504 3803 524
rect 3811 504 3823 584
rect 3842 504 3854 584
rect 3870 504 3882 584
rect 3892 504 3904 544
rect 3951 504 3963 544
rect 3971 504 3983 544
rect 3991 504 4003 544
rect 4017 504 4029 584
rect 4037 504 4049 524
rect 4067 504 4079 524
rect 4095 504 4107 544
rect 4121 504 4133 544
rect 4141 504 4153 544
rect 4173 504 4185 544
rect 4207 504 4219 544
rect 4227 504 4239 584
rect 4257 504 4269 544
rect 4277 504 4289 544
rect 4297 504 4309 544
rect 4337 504 4349 544
rect 4357 504 4369 544
rect 4377 504 4389 544
rect 4436 504 4448 544
rect 4458 504 4470 584
rect 4486 504 4498 584
rect 4521 504 4533 584
rect 4541 504 4553 544
rect 4575 504 4587 544
rect 4607 504 4619 544
rect 4627 504 4639 544
rect 4653 504 4665 544
rect 4681 504 4693 524
rect 4711 504 4723 524
rect 4731 504 4743 584
rect 17 436 29 476
rect 37 436 49 476
rect 57 436 69 476
rect 97 436 109 476
rect 117 436 129 476
rect 137 436 149 476
rect 191 436 203 476
rect 211 436 223 476
rect 231 436 243 476
rect 271 436 283 476
rect 291 436 303 476
rect 311 436 323 476
rect 347 396 359 476
rect 367 396 379 476
rect 391 436 403 476
rect 411 436 423 476
rect 451 436 463 476
rect 471 436 483 476
rect 491 436 503 476
rect 531 436 543 476
rect 551 440 563 476
rect 571 436 583 476
rect 591 436 603 476
rect 631 396 643 476
rect 651 396 663 464
rect 671 398 683 476
rect 691 410 703 476
rect 711 398 723 476
rect 763 396 775 476
rect 791 396 803 476
rect 831 436 843 476
rect 851 436 863 476
rect 871 436 883 476
rect 897 436 909 476
rect 917 436 929 476
rect 937 436 949 476
rect 991 436 1003 476
rect 1011 436 1023 476
rect 1031 436 1043 476
rect 1071 436 1083 476
rect 1091 436 1103 476
rect 1111 436 1123 476
rect 1151 396 1163 476
rect 1171 396 1183 464
rect 1191 398 1203 476
rect 1211 410 1223 476
rect 1231 398 1243 476
rect 1262 396 1274 476
rect 1290 396 1302 476
rect 1312 436 1324 476
rect 1383 396 1395 476
rect 1411 396 1423 476
rect 1442 396 1454 476
rect 1470 396 1482 476
rect 1492 436 1504 476
rect 1537 436 1549 476
rect 1557 436 1569 476
rect 1611 396 1623 476
rect 1631 396 1643 476
rect 1651 408 1663 476
rect 1671 404 1683 476
rect 1697 436 1709 476
rect 1717 436 1729 476
rect 1757 436 1769 476
rect 1777 436 1789 476
rect 1797 440 1809 476
rect 1817 436 1829 476
rect 1857 404 1869 476
rect 1877 408 1889 476
rect 1897 396 1909 476
rect 1917 396 1929 476
rect 1957 436 1969 476
rect 1977 436 1989 476
rect 1997 436 2009 476
rect 2037 436 2049 476
rect 2057 436 2069 476
rect 2077 436 2089 476
rect 2117 436 2129 476
rect 2137 436 2149 476
rect 2157 436 2169 476
rect 2223 396 2235 476
rect 2251 396 2263 476
rect 2291 436 2303 476
rect 2311 436 2323 476
rect 2331 436 2343 476
rect 2357 396 2369 476
rect 2385 396 2397 476
rect 2437 436 2449 476
rect 2457 436 2469 476
rect 2477 440 2489 476
rect 2497 436 2509 476
rect 2551 436 2563 476
rect 2571 436 2583 476
rect 2611 436 2623 476
rect 2631 440 2643 476
rect 2651 436 2663 476
rect 2671 436 2683 476
rect 2697 404 2709 476
rect 2717 408 2729 476
rect 2737 396 2749 476
rect 2757 396 2769 476
rect 2797 396 2809 476
rect 2825 396 2837 476
rect 2891 436 2903 476
rect 2911 436 2923 476
rect 2931 436 2943 476
rect 2976 436 2988 476
rect 2998 396 3010 476
rect 3026 396 3038 476
rect 3076 436 3088 476
rect 3098 396 3110 476
rect 3126 396 3138 476
rect 3183 396 3195 476
rect 3211 396 3223 476
rect 3251 436 3263 476
rect 3271 436 3283 476
rect 3316 436 3328 476
rect 3338 396 3350 476
rect 3366 396 3378 476
rect 3411 396 3423 476
rect 3431 396 3443 476
rect 3451 408 3463 476
rect 3471 404 3483 476
rect 3523 396 3535 476
rect 3551 396 3563 476
rect 3577 396 3589 476
rect 3607 397 3619 476
rect 3627 397 3639 476
rect 3677 436 3689 476
rect 3697 436 3709 476
rect 3717 436 3729 476
rect 3757 436 3769 476
rect 3777 436 3789 476
rect 3797 436 3809 476
rect 3856 436 3868 476
rect 3878 396 3890 476
rect 3906 396 3918 476
rect 3951 436 3963 476
rect 3971 436 3983 476
rect 4011 436 4023 476
rect 4031 436 4043 476
rect 4057 396 4069 476
rect 4077 456 4089 476
rect 4107 456 4119 476
rect 4135 436 4147 476
rect 4161 436 4173 476
rect 4181 436 4193 476
rect 4213 436 4225 476
rect 4247 436 4259 476
rect 4267 396 4279 476
rect 4311 436 4323 476
rect 4331 436 4343 476
rect 4351 436 4363 476
rect 4396 436 4408 476
rect 4418 396 4430 476
rect 4446 396 4458 476
rect 4491 436 4503 476
rect 4511 436 4523 476
rect 4537 396 4549 476
rect 4557 456 4569 476
rect 4587 456 4599 476
rect 4615 436 4627 476
rect 4641 436 4653 476
rect 4661 436 4673 476
rect 4693 436 4705 476
rect 4727 436 4739 476
rect 4747 396 4759 476
rect 31 24 43 64
rect 51 24 63 60
rect 71 24 83 64
rect 91 24 103 64
rect 117 24 129 96
rect 137 24 149 92
rect 157 24 169 104
rect 177 24 189 104
rect 236 24 248 64
rect 258 24 270 104
rect 286 24 298 104
rect 322 24 334 104
rect 350 24 362 104
rect 372 24 384 64
rect 431 24 443 64
rect 451 24 463 60
rect 471 24 483 64
rect 491 24 503 64
rect 517 24 529 64
rect 537 24 549 64
rect 557 24 569 60
rect 577 24 589 64
rect 617 24 629 96
rect 637 24 649 92
rect 657 24 669 104
rect 677 24 689 104
rect 731 24 743 104
rect 751 24 763 104
rect 771 24 783 92
rect 791 24 803 96
rect 817 24 829 64
rect 837 24 849 64
rect 896 24 908 64
rect 918 24 930 104
rect 946 24 958 104
rect 991 24 1003 64
rect 1011 24 1023 64
rect 1042 24 1054 104
rect 1070 24 1082 104
rect 1092 24 1104 64
rect 1142 24 1154 104
rect 1170 24 1182 104
rect 1192 24 1204 64
rect 1237 24 1249 64
rect 1257 24 1269 64
rect 1277 24 1289 60
rect 1297 24 1309 64
rect 1337 24 1349 64
rect 1357 24 1369 64
rect 1377 24 1389 60
rect 1397 24 1409 64
rect 1451 24 1463 104
rect 1471 24 1483 104
rect 1491 24 1503 92
rect 1511 24 1523 96
rect 1537 24 1549 64
rect 1557 24 1569 64
rect 1577 24 1589 60
rect 1597 24 1609 64
rect 1651 24 1663 104
rect 1671 24 1683 104
rect 1691 24 1703 92
rect 1711 24 1723 96
rect 1737 24 1749 64
rect 1757 24 1769 64
rect 1777 24 1789 60
rect 1797 24 1809 64
rect 1837 24 1849 64
rect 1857 24 1869 64
rect 1877 24 1889 64
rect 1917 24 1929 64
rect 1939 24 1951 104
rect 1959 24 1971 104
rect 2007 24 2019 104
rect 2027 24 2039 104
rect 2051 24 2063 64
rect 2071 24 2083 64
rect 2097 24 2109 64
rect 2119 24 2131 104
rect 2139 24 2151 104
rect 2177 24 2189 64
rect 2197 24 2209 64
rect 2217 24 2229 60
rect 2237 24 2249 64
rect 2277 24 2289 102
rect 2297 24 2309 90
rect 2317 24 2329 102
rect 2337 36 2349 104
rect 2357 24 2369 104
rect 2402 24 2414 104
rect 2430 24 2442 104
rect 2452 24 2464 64
rect 2511 24 2523 104
rect 2531 24 2543 104
rect 2551 24 2563 92
rect 2571 24 2583 96
rect 2602 24 2614 104
rect 2630 24 2642 104
rect 2652 24 2664 64
rect 2697 24 2709 64
rect 2717 24 2729 64
rect 2757 24 2769 64
rect 2777 24 2789 64
rect 2797 24 2809 60
rect 2817 24 2829 64
rect 2857 24 2869 64
rect 2877 24 2889 64
rect 2921 24 2933 104
rect 2941 24 2953 64
rect 2975 24 2987 64
rect 3007 24 3019 64
rect 3027 24 3039 64
rect 3053 24 3065 64
rect 3081 24 3093 44
rect 3111 24 3123 44
rect 3131 24 3143 104
rect 3157 24 3169 64
rect 3177 24 3189 64
rect 3231 24 3243 64
rect 3251 24 3263 64
rect 3281 24 3293 104
rect 3301 24 3313 64
rect 3335 24 3347 64
rect 3367 24 3379 64
rect 3387 24 3399 64
rect 3413 24 3425 64
rect 3441 24 3453 44
rect 3471 24 3483 44
rect 3491 24 3503 104
rect 3543 24 3555 104
rect 3571 24 3583 104
rect 3597 24 3609 104
rect 3617 24 3629 44
rect 3647 24 3659 44
rect 3675 24 3687 64
rect 3701 24 3713 64
rect 3721 24 3733 64
rect 3753 24 3765 64
rect 3787 24 3799 64
rect 3807 24 3819 104
rect 3837 24 3849 64
rect 3857 24 3869 64
rect 3902 24 3914 104
rect 3930 24 3942 104
rect 3952 24 3964 64
rect 3997 24 4009 104
rect 4025 24 4037 104
rect 4077 24 4089 104
rect 4105 24 4117 104
rect 4183 24 4195 104
rect 4211 24 4223 104
rect 4242 24 4254 104
rect 4270 24 4282 104
rect 4292 24 4304 64
rect 4351 24 4363 64
rect 4371 24 4383 64
rect 4391 24 4403 64
rect 4431 24 4443 64
rect 4451 24 4463 64
rect 4477 24 4489 104
rect 4505 24 4517 104
rect 4557 24 4569 64
rect 4577 24 4589 64
rect 4597 24 4609 64
rect 4651 24 4663 64
rect 4671 24 4683 64
rect 4697 24 4709 64
rect 4717 24 4729 64
rect 4737 24 4749 64
<< psubstratepcontact >>
rect 4 4564 4776 4576
rect 4 4084 4776 4096
rect 4 3604 4776 3616
rect 4 3124 4776 3136
rect 4 2644 4776 2656
rect 4 2164 4776 2176
rect 4 1684 4776 1696
rect 4 1204 4776 1216
rect 4 724 4776 736
rect 4 244 4776 256
<< nsubstratencontact >>
rect 4 4324 4776 4336
rect 4 3844 4776 3856
rect 4 3364 4776 3376
rect 4 2884 4776 2896
rect 4 2404 4776 2416
rect 4 1924 4776 1936
rect 4 1444 4776 1456
rect 4 964 4776 976
rect 4 484 4776 496
rect 4 4 4776 16
<< polysilicon >>
rect 52 4556 56 4560
rect 74 4556 78 4560
rect 82 4556 86 4560
rect 168 4556 172 4560
rect 176 4556 180 4560
rect 184 4556 188 4560
rect 232 4556 236 4560
rect 240 4556 244 4560
rect 248 4556 252 4560
rect 368 4556 372 4560
rect 376 4556 380 4560
rect 384 4556 388 4560
rect 434 4556 438 4560
rect 442 4556 446 4560
rect 464 4556 468 4560
rect 531 4556 535 4560
rect 551 4556 555 4560
rect 571 4556 575 4560
rect 631 4556 635 4560
rect 651 4556 655 4560
rect 671 4556 675 4560
rect 768 4556 772 4560
rect 776 4556 780 4560
rect 784 4556 788 4560
rect 832 4556 836 4560
rect 840 4556 844 4560
rect 848 4556 852 4560
rect 933 4556 937 4560
rect 943 4556 947 4560
rect 1012 4556 1016 4560
rect 1020 4556 1024 4560
rect 1028 4556 1032 4560
rect 1114 4556 1118 4560
rect 1122 4556 1126 4560
rect 1144 4556 1148 4560
rect 1233 4556 1237 4560
rect 1243 4556 1247 4560
rect 1305 4556 1309 4560
rect 1325 4556 1329 4560
rect 1385 4556 1389 4560
rect 1405 4556 1409 4560
rect 1425 4556 1429 4560
rect 1493 4556 1497 4560
rect 1503 4556 1507 4560
rect 1551 4556 1555 4560
rect 1571 4556 1575 4560
rect 1632 4556 1636 4560
rect 1640 4556 1644 4560
rect 1648 4556 1652 4560
rect 1752 4556 1756 4560
rect 1774 4556 1778 4560
rect 1782 4556 1786 4560
rect 1831 4556 1835 4560
rect 1905 4556 1909 4560
rect 1954 4556 1958 4560
rect 1962 4556 1966 4560
rect 1984 4556 1988 4560
rect 2051 4556 2055 4560
rect 2071 4556 2075 4560
rect 2131 4556 2135 4560
rect 2191 4556 2195 4560
rect 2211 4556 2215 4560
rect 2231 4556 2235 4560
rect 2305 4556 2309 4560
rect 2325 4556 2329 4560
rect 2345 4556 2349 4560
rect 2365 4556 2369 4560
rect 2411 4556 2415 4560
rect 2431 4556 2435 4560
rect 2451 4556 2455 4560
rect 2514 4556 2518 4560
rect 2522 4556 2526 4560
rect 2544 4556 2548 4560
rect 2646 4556 2650 4560
rect 2654 4556 2658 4560
rect 2674 4556 2678 4560
rect 2682 4556 2686 4560
rect 2735 4556 2739 4560
rect 2755 4556 2759 4560
rect 2765 4556 2769 4560
rect 2787 4556 2791 4560
rect 2797 4556 2801 4560
rect 2819 4556 2823 4560
rect 2865 4556 2869 4560
rect 2873 4556 2877 4560
rect 2893 4556 2897 4560
rect 2903 4556 2907 4560
rect 2925 4556 2929 4560
rect 2985 4556 2989 4560
rect 3045 4556 3049 4560
rect 3065 4556 3069 4560
rect 3085 4556 3089 4560
rect 3145 4556 3149 4560
rect 3165 4556 3169 4560
rect 3225 4556 3229 4560
rect 3245 4556 3249 4560
rect 3265 4556 3269 4560
rect 3325 4556 3329 4560
rect 3345 4556 3349 4560
rect 3405 4556 3409 4560
rect 3451 4556 3455 4560
rect 3473 4556 3477 4560
rect 3483 4556 3487 4560
rect 3503 4556 3507 4560
rect 3511 4556 3515 4560
rect 3557 4556 3561 4560
rect 3579 4556 3583 4560
rect 3589 4556 3593 4560
rect 3611 4556 3615 4560
rect 3621 4556 3625 4560
rect 3641 4556 3645 4560
rect 3691 4556 3695 4560
rect 3711 4556 3715 4560
rect 3731 4556 3735 4560
rect 3793 4556 3797 4560
rect 3803 4556 3807 4560
rect 3885 4556 3889 4560
rect 3905 4556 3909 4560
rect 3925 4556 3929 4560
rect 3945 4556 3949 4560
rect 3965 4556 3969 4560
rect 3985 4556 3989 4560
rect 4005 4556 4009 4560
rect 4025 4556 4029 4560
rect 4083 4556 4087 4560
rect 4105 4556 4109 4560
rect 4153 4556 4157 4560
rect 4163 4556 4167 4560
rect 4231 4556 4235 4560
rect 4291 4556 4295 4560
rect 4311 4556 4315 4560
rect 4331 4556 4335 4560
rect 4391 4556 4395 4560
rect 4413 4556 4417 4560
rect 4423 4556 4427 4560
rect 4443 4556 4447 4560
rect 4451 4556 4455 4560
rect 4497 4556 4501 4560
rect 4519 4556 4523 4560
rect 4529 4556 4533 4560
rect 4551 4556 4555 4560
rect 4561 4556 4565 4560
rect 4581 4556 4585 4560
rect 4631 4556 4635 4560
rect 4653 4556 4657 4560
rect 4713 4556 4717 4560
rect 4723 4556 4727 4560
rect 52 4493 56 4536
rect 45 4481 54 4493
rect 45 4424 49 4481
rect 74 4479 78 4516
rect 82 4512 86 4516
rect 82 4506 101 4512
rect 94 4493 101 4506
rect 434 4512 438 4516
rect 419 4506 438 4512
rect 74 4444 80 4467
rect 94 4444 101 4481
rect 65 4438 80 4444
rect 85 4438 101 4444
rect 168 4439 172 4496
rect 65 4424 69 4438
rect 85 4424 89 4438
rect 145 4427 153 4439
rect 165 4427 172 4439
rect 145 4384 149 4427
rect 176 4419 180 4496
rect 184 4439 188 4496
rect 232 4439 236 4496
rect 184 4427 194 4439
rect 226 4427 236 4439
rect 174 4400 180 4407
rect 165 4396 180 4400
rect 194 4396 200 4427
rect 165 4384 169 4396
rect 185 4392 200 4396
rect 220 4396 226 4427
rect 240 4419 244 4496
rect 248 4439 252 4496
rect 368 4439 372 4496
rect 248 4427 255 4439
rect 267 4427 275 4439
rect 240 4400 246 4407
rect 240 4396 255 4400
rect 220 4392 235 4396
rect 185 4384 189 4392
rect 231 4384 235 4392
rect 251 4384 255 4396
rect 271 4384 275 4427
rect 345 4427 353 4439
rect 365 4427 372 4439
rect 345 4384 349 4427
rect 376 4419 380 4496
rect 384 4439 388 4496
rect 419 4493 426 4506
rect 419 4444 426 4481
rect 442 4479 446 4516
rect 464 4493 468 4536
rect 531 4511 535 4516
rect 522 4504 535 4511
rect 466 4481 475 4493
rect 440 4444 446 4467
rect 384 4427 394 4439
rect 419 4438 435 4444
rect 440 4438 455 4444
rect 374 4400 380 4407
rect 365 4396 380 4400
rect 394 4396 400 4427
rect 431 4424 435 4438
rect 451 4424 455 4438
rect 471 4424 475 4481
rect 522 4459 526 4504
rect 551 4493 555 4516
rect 546 4481 555 4493
rect 522 4436 526 4447
rect 522 4428 540 4436
rect 536 4424 540 4428
rect 544 4424 548 4481
rect 571 4439 575 4516
rect 631 4511 635 4516
rect 622 4504 635 4511
rect 622 4459 626 4504
rect 651 4493 655 4516
rect 646 4481 655 4493
rect 566 4427 573 4439
rect 622 4436 626 4447
rect 622 4428 640 4436
rect 365 4384 369 4396
rect 385 4392 400 4396
rect 385 4384 389 4392
rect 566 4384 570 4427
rect 636 4424 640 4428
rect 644 4424 648 4481
rect 671 4439 675 4516
rect 933 4496 937 4516
rect 768 4439 772 4496
rect 666 4427 673 4439
rect 745 4427 753 4439
rect 765 4427 772 4439
rect 666 4384 670 4427
rect 745 4384 749 4427
rect 776 4419 780 4496
rect 784 4439 788 4496
rect 832 4439 836 4496
rect 784 4427 794 4439
rect 826 4427 836 4439
rect 774 4400 780 4407
rect 765 4396 780 4400
rect 794 4396 800 4427
rect 765 4384 769 4396
rect 785 4392 800 4396
rect 820 4396 826 4427
rect 840 4419 844 4496
rect 848 4439 852 4496
rect 929 4489 937 4496
rect 943 4496 947 4516
rect 1114 4512 1118 4516
rect 1099 4506 1118 4512
rect 943 4489 957 4496
rect 929 4473 935 4489
rect 926 4461 935 4473
rect 848 4427 855 4439
rect 867 4427 875 4439
rect 840 4400 846 4407
rect 840 4396 855 4400
rect 820 4392 835 4396
rect 785 4384 789 4392
rect 831 4384 835 4392
rect 851 4384 855 4396
rect 871 4384 875 4427
rect 931 4384 935 4461
rect 951 4473 957 4489
rect 951 4461 954 4473
rect 951 4384 955 4461
rect 1012 4439 1016 4496
rect 1006 4427 1016 4439
rect 1000 4396 1006 4427
rect 1020 4419 1024 4496
rect 1028 4439 1032 4496
rect 1099 4493 1106 4506
rect 1099 4444 1106 4481
rect 1122 4479 1126 4516
rect 1144 4493 1148 4536
rect 1233 4496 1237 4516
rect 1146 4481 1155 4493
rect 1120 4444 1126 4467
rect 1028 4427 1035 4439
rect 1047 4427 1055 4439
rect 1099 4438 1115 4444
rect 1120 4438 1135 4444
rect 1020 4400 1026 4407
rect 1020 4396 1035 4400
rect 1000 4392 1015 4396
rect 1011 4384 1015 4392
rect 1031 4384 1035 4396
rect 1051 4384 1055 4427
rect 1111 4424 1115 4438
rect 1131 4424 1135 4438
rect 1151 4424 1155 4481
rect 1223 4489 1237 4496
rect 1243 4496 1247 4516
rect 1243 4489 1251 4496
rect 1223 4473 1229 4489
rect 1226 4461 1229 4473
rect 1225 4384 1229 4461
rect 1245 4473 1251 4489
rect 1245 4461 1254 4473
rect 1245 4384 1249 4461
rect 1305 4459 1309 4536
rect 1325 4459 1329 4536
rect 1306 4447 1321 4459
rect 1317 4424 1321 4447
rect 1325 4447 1334 4459
rect 1325 4424 1329 4447
rect 1385 4439 1389 4516
rect 1405 4493 1409 4516
rect 1425 4511 1429 4516
rect 1425 4504 1438 4511
rect 1405 4481 1414 4493
rect 1387 4427 1394 4439
rect 1390 4384 1394 4427
rect 1412 4424 1416 4481
rect 1434 4459 1438 4504
rect 1493 4496 1497 4516
rect 1483 4489 1497 4496
rect 1503 4496 1507 4516
rect 1503 4489 1511 4496
rect 1483 4473 1489 4489
rect 1486 4461 1489 4473
rect 1434 4436 1438 4447
rect 1420 4428 1438 4436
rect 1420 4424 1424 4428
rect 1485 4384 1489 4461
rect 1505 4473 1511 4489
rect 1505 4461 1514 4473
rect 1505 4384 1509 4461
rect 1551 4459 1555 4536
rect 1571 4459 1575 4536
rect 1546 4447 1555 4459
rect 1551 4424 1555 4447
rect 1559 4447 1574 4459
rect 1559 4424 1563 4447
rect 1632 4439 1636 4496
rect 1626 4427 1636 4439
rect 1620 4396 1626 4427
rect 1640 4419 1644 4496
rect 1648 4439 1652 4496
rect 1752 4493 1756 4536
rect 1745 4481 1754 4493
rect 1648 4427 1655 4439
rect 1667 4427 1675 4439
rect 1640 4400 1646 4407
rect 1640 4396 1655 4400
rect 1620 4392 1635 4396
rect 1631 4384 1635 4392
rect 1651 4384 1655 4396
rect 1671 4384 1675 4427
rect 1745 4424 1749 4481
rect 1774 4479 1778 4516
rect 1782 4512 1786 4516
rect 1782 4506 1801 4512
rect 1794 4493 1801 4506
rect 1774 4444 1780 4467
rect 1794 4444 1801 4481
rect 1831 4479 1835 4536
rect 1826 4467 1835 4479
rect 1765 4438 1780 4444
rect 1785 4438 1801 4444
rect 1765 4424 1769 4438
rect 1785 4424 1789 4438
rect 1831 4384 1835 4467
rect 1905 4479 1909 4536
rect 1954 4512 1958 4516
rect 1939 4506 1958 4512
rect 1939 4493 1946 4506
rect 1905 4467 1914 4479
rect 1905 4384 1909 4467
rect 1939 4444 1946 4481
rect 1962 4479 1966 4516
rect 1984 4493 1988 4536
rect 1986 4481 1995 4493
rect 1960 4444 1966 4467
rect 1939 4438 1955 4444
rect 1960 4438 1975 4444
rect 1951 4424 1955 4438
rect 1971 4424 1975 4438
rect 1991 4424 1995 4481
rect 2051 4459 2055 4536
rect 2071 4459 2075 4536
rect 2131 4479 2135 4536
rect 2411 4529 2415 4536
rect 2431 4529 2435 4536
rect 2402 4524 2415 4529
rect 2191 4511 2195 4516
rect 2126 4467 2135 4479
rect 2046 4447 2055 4459
rect 2051 4424 2055 4447
rect 2059 4447 2074 4459
rect 2059 4424 2063 4447
rect 2131 4384 2135 4467
rect 2182 4504 2195 4511
rect 2182 4459 2186 4504
rect 2211 4493 2215 4516
rect 2206 4481 2215 4493
rect 2182 4436 2186 4447
rect 2182 4428 2200 4436
rect 2196 4424 2200 4428
rect 2204 4424 2208 4481
rect 2231 4439 2235 4516
rect 2305 4459 2309 4516
rect 2325 4493 2329 4516
rect 2345 4493 2349 4516
rect 2365 4509 2369 4516
rect 2365 4505 2380 4509
rect 2345 4481 2354 4493
rect 2307 4447 2309 4459
rect 2226 4427 2233 4439
rect 2305 4432 2309 4447
rect 2305 4428 2319 4432
rect 2226 4384 2230 4427
rect 2315 4424 2319 4428
rect 2325 4424 2329 4481
rect 2345 4432 2351 4481
rect 2374 4459 2380 4505
rect 2402 4479 2406 4524
rect 2374 4432 2379 4447
rect 2345 4428 2359 4432
rect 2355 4424 2359 4428
rect 2365 4428 2379 4432
rect 2402 4433 2406 4467
rect 2421 4523 2435 4529
rect 2421 4459 2425 4523
rect 2451 4508 2455 4516
rect 2514 4512 2518 4516
rect 2445 4496 2455 4508
rect 2499 4506 2518 4512
rect 2499 4493 2506 4506
rect 2402 4428 2415 4433
rect 2365 4424 2369 4428
rect 2411 4424 2415 4428
rect 2421 4424 2425 4447
rect 2499 4444 2506 4481
rect 2522 4479 2526 4516
rect 2544 4493 2548 4536
rect 2646 4511 2650 4516
rect 2620 4507 2650 4511
rect 2546 4481 2555 4493
rect 2520 4444 2526 4467
rect 2499 4438 2515 4444
rect 2520 4438 2535 4444
rect 2441 4424 2445 4429
rect 2511 4424 2515 4438
rect 2531 4424 2535 4438
rect 2551 4424 2555 4481
rect 2620 4459 2626 4507
rect 2654 4502 2658 4516
rect 2645 4495 2658 4502
rect 2645 4493 2649 4495
rect 2674 4493 2678 4516
rect 2682 4508 2686 4516
rect 2682 4501 2699 4508
rect 2647 4481 2649 4493
rect 2626 4447 2629 4459
rect 2625 4424 2629 4447
rect 2645 4424 2649 4481
rect 2674 4452 2678 4481
rect 2693 4459 2699 4501
rect 2735 4479 2739 4516
rect 2755 4478 2759 4536
rect 2765 4504 2769 4536
rect 2787 4524 2791 4536
rect 2789 4512 2791 4524
rect 2797 4524 2801 4536
rect 2797 4512 2799 4524
rect 2765 4500 2798 4504
rect 2665 4446 2678 4452
rect 2685 4447 2693 4452
rect 2685 4446 2705 4447
rect 2665 4424 2669 4446
rect 2685 4424 2689 4446
rect 2735 4424 2739 4467
rect 2755 4384 2759 4466
rect 2774 4451 2778 4480
rect 2769 4443 2778 4451
rect 2769 4384 2773 4443
rect 2794 4436 2798 4500
rect 2795 4424 2798 4436
rect 2789 4384 2793 4424
rect 2803 4402 2807 4512
rect 2819 4422 2823 4536
rect 2865 4532 2869 4536
rect 2835 4528 2869 4532
rect 2801 4384 2805 4390
rect 2821 4384 2825 4410
rect 2835 4402 2839 4528
rect 2873 4524 2877 4536
rect 2847 4520 2877 4524
rect 2859 4519 2877 4520
rect 2893 4515 2897 4536
rect 2873 4511 2897 4515
rect 2873 4416 2879 4511
rect 2903 4487 2907 4536
rect 2903 4429 2907 4475
rect 2925 4448 2929 4516
rect 2927 4436 2929 4448
rect 2903 4423 2911 4429
rect 2925 4424 2929 4436
rect 2985 4479 2989 4536
rect 2985 4467 2994 4479
rect 2847 4390 2871 4392
rect 2835 4388 2871 4390
rect 2867 4384 2871 4388
rect 2875 4384 2879 4416
rect 2895 4364 2899 4404
rect 2907 4394 2911 4423
rect 2903 4387 2911 4394
rect 2903 4364 2907 4387
rect 2985 4384 2989 4467
rect 3045 4439 3049 4516
rect 3065 4493 3069 4516
rect 3085 4511 3089 4516
rect 3085 4504 3098 4511
rect 3065 4481 3074 4493
rect 3047 4427 3054 4439
rect 3050 4384 3054 4427
rect 3072 4424 3076 4481
rect 3094 4459 3098 4504
rect 3145 4459 3149 4536
rect 3165 4459 3169 4536
rect 3146 4447 3161 4459
rect 3094 4436 3098 4447
rect 3080 4428 3098 4436
rect 3080 4424 3084 4428
rect 3157 4424 3161 4447
rect 3165 4447 3174 4459
rect 3165 4424 3169 4447
rect 3225 4439 3229 4516
rect 3245 4493 3249 4516
rect 3265 4511 3269 4516
rect 3265 4504 3278 4511
rect 3245 4481 3254 4493
rect 3227 4427 3234 4439
rect 3230 4384 3234 4427
rect 3252 4424 3256 4481
rect 3274 4459 3278 4504
rect 3325 4459 3329 4536
rect 3345 4459 3349 4536
rect 3405 4479 3409 4536
rect 3405 4467 3414 4479
rect 3326 4447 3341 4459
rect 3274 4436 3278 4447
rect 3260 4428 3278 4436
rect 3260 4424 3264 4428
rect 3337 4424 3341 4447
rect 3345 4447 3354 4459
rect 3345 4424 3349 4447
rect 3405 4384 3409 4467
rect 3451 4448 3455 4516
rect 3473 4487 3477 4536
rect 3483 4515 3487 4536
rect 3503 4524 3507 4536
rect 3511 4532 3515 4536
rect 3511 4528 3545 4532
rect 3503 4520 3533 4524
rect 3503 4519 3521 4520
rect 3483 4511 3507 4515
rect 3451 4436 3453 4448
rect 3451 4424 3455 4436
rect 3473 4429 3477 4475
rect 3469 4423 3477 4429
rect 3469 4394 3473 4423
rect 3501 4416 3507 4511
rect 3469 4387 3477 4394
rect 3473 4364 3477 4387
rect 3481 4364 3485 4404
rect 3501 4384 3505 4416
rect 3541 4402 3545 4528
rect 3557 4422 3561 4536
rect 3579 4524 3583 4536
rect 3581 4512 3583 4524
rect 3589 4524 3593 4536
rect 3589 4512 3591 4524
rect 3509 4390 3533 4392
rect 3509 4388 3545 4390
rect 3509 4384 3513 4388
rect 3555 4384 3559 4410
rect 3573 4402 3577 4512
rect 3611 4504 3615 4536
rect 3582 4500 3615 4504
rect 3582 4436 3586 4500
rect 3602 4451 3606 4480
rect 3621 4478 3625 4536
rect 3641 4479 3645 4516
rect 3691 4511 3695 4516
rect 3682 4504 3695 4511
rect 3602 4443 3611 4451
rect 3582 4424 3585 4436
rect 3575 4384 3579 4390
rect 3587 4384 3591 4424
rect 3607 4384 3611 4443
rect 3621 4384 3625 4466
rect 3641 4424 3645 4467
rect 3682 4459 3686 4504
rect 3711 4493 3715 4516
rect 3706 4481 3715 4493
rect 3682 4436 3686 4447
rect 3682 4428 3700 4436
rect 3696 4424 3700 4428
rect 3704 4424 3708 4481
rect 3731 4439 3735 4516
rect 3793 4496 3797 4516
rect 3789 4489 3797 4496
rect 3803 4496 3807 4516
rect 3885 4496 3889 4516
rect 3905 4496 3909 4516
rect 3925 4496 3929 4516
rect 3945 4496 3949 4516
rect 3965 4496 3969 4516
rect 3985 4496 3989 4516
rect 3803 4489 3817 4496
rect 3789 4473 3795 4489
rect 3786 4461 3795 4473
rect 3726 4427 3733 4439
rect 3726 4384 3730 4427
rect 3791 4384 3795 4461
rect 3811 4473 3817 4489
rect 3885 4484 3898 4496
rect 3925 4484 3938 4496
rect 3965 4484 3978 4496
rect 4005 4493 4009 4516
rect 4025 4493 4029 4516
rect 4083 4510 4087 4516
rect 4083 4498 4085 4510
rect 3811 4461 3814 4473
rect 3811 4384 3815 4461
rect 3885 4424 3889 4484
rect 3905 4424 3909 4484
rect 3925 4424 3929 4484
rect 3945 4424 3949 4484
rect 3965 4424 3969 4484
rect 3985 4424 3989 4484
rect 4005 4481 4014 4493
rect 4026 4481 4029 4493
rect 4005 4424 4009 4481
rect 4025 4424 4029 4481
rect 4105 4459 4109 4536
rect 4153 4496 4157 4516
rect 4149 4489 4157 4496
rect 4163 4496 4167 4516
rect 4163 4489 4177 4496
rect 4149 4473 4155 4489
rect 4146 4461 4155 4473
rect 4105 4447 4114 4459
rect 4083 4430 4085 4442
rect 4083 4424 4087 4430
rect 4105 4384 4109 4447
rect 4151 4384 4155 4461
rect 4171 4473 4177 4489
rect 4231 4479 4235 4536
rect 4291 4511 4295 4516
rect 4171 4461 4174 4473
rect 4226 4467 4235 4479
rect 4171 4384 4175 4461
rect 4231 4384 4235 4467
rect 4282 4504 4295 4511
rect 4282 4459 4286 4504
rect 4311 4493 4315 4516
rect 4306 4481 4315 4493
rect 4282 4436 4286 4447
rect 4282 4428 4300 4436
rect 4296 4424 4300 4428
rect 4304 4424 4308 4481
rect 4331 4439 4335 4516
rect 4391 4448 4395 4516
rect 4413 4487 4417 4536
rect 4423 4515 4427 4536
rect 4443 4524 4447 4536
rect 4451 4532 4455 4536
rect 4451 4528 4485 4532
rect 4443 4520 4473 4524
rect 4443 4519 4461 4520
rect 4423 4511 4447 4515
rect 4326 4427 4333 4439
rect 4391 4436 4393 4448
rect 4326 4384 4330 4427
rect 4391 4424 4395 4436
rect 4413 4429 4417 4475
rect 4409 4423 4417 4429
rect 4409 4394 4413 4423
rect 4441 4416 4447 4511
rect 4409 4387 4417 4394
rect 4413 4364 4417 4387
rect 4421 4364 4425 4404
rect 4441 4384 4445 4416
rect 4481 4402 4485 4528
rect 4497 4422 4501 4536
rect 4519 4524 4523 4536
rect 4521 4512 4523 4524
rect 4529 4524 4533 4536
rect 4529 4512 4531 4524
rect 4449 4390 4473 4392
rect 4449 4388 4485 4390
rect 4449 4384 4453 4388
rect 4495 4384 4499 4410
rect 4513 4402 4517 4512
rect 4551 4504 4555 4536
rect 4522 4500 4555 4504
rect 4522 4436 4526 4500
rect 4542 4451 4546 4480
rect 4561 4478 4565 4536
rect 4581 4479 4585 4516
rect 4542 4443 4551 4451
rect 4522 4424 4525 4436
rect 4515 4384 4519 4390
rect 4527 4384 4531 4424
rect 4547 4384 4551 4443
rect 4561 4384 4565 4466
rect 4581 4424 4585 4467
rect 4631 4459 4635 4536
rect 4653 4510 4657 4516
rect 4655 4498 4657 4510
rect 4713 4496 4717 4516
rect 4709 4489 4717 4496
rect 4723 4496 4727 4516
rect 4723 4489 4737 4496
rect 4709 4473 4715 4489
rect 4706 4461 4715 4473
rect 4626 4447 4635 4459
rect 4631 4384 4635 4447
rect 4655 4430 4657 4442
rect 4653 4424 4657 4430
rect 4711 4384 4715 4461
rect 4731 4473 4737 4489
rect 4731 4461 4734 4473
rect 4731 4384 4735 4461
rect 45 4340 49 4344
rect 65 4340 69 4344
rect 85 4340 89 4344
rect 145 4340 149 4344
rect 165 4340 169 4344
rect 185 4340 189 4344
rect 231 4340 235 4344
rect 251 4340 255 4344
rect 271 4340 275 4344
rect 345 4340 349 4344
rect 365 4340 369 4344
rect 385 4340 389 4344
rect 431 4340 435 4344
rect 451 4340 455 4344
rect 471 4340 475 4344
rect 536 4340 540 4344
rect 544 4340 548 4344
rect 566 4340 570 4344
rect 636 4340 640 4344
rect 644 4340 648 4344
rect 666 4340 670 4344
rect 745 4340 749 4344
rect 765 4340 769 4344
rect 785 4340 789 4344
rect 831 4340 835 4344
rect 851 4340 855 4344
rect 871 4340 875 4344
rect 931 4340 935 4344
rect 951 4340 955 4344
rect 1011 4340 1015 4344
rect 1031 4340 1035 4344
rect 1051 4340 1055 4344
rect 1111 4340 1115 4344
rect 1131 4340 1135 4344
rect 1151 4340 1155 4344
rect 1225 4340 1229 4344
rect 1245 4340 1249 4344
rect 1317 4340 1321 4344
rect 1325 4340 1329 4344
rect 1390 4340 1394 4344
rect 1412 4340 1416 4344
rect 1420 4340 1424 4344
rect 1485 4340 1489 4344
rect 1505 4340 1509 4344
rect 1551 4340 1555 4344
rect 1559 4340 1563 4344
rect 1631 4340 1635 4344
rect 1651 4340 1655 4344
rect 1671 4340 1675 4344
rect 1745 4340 1749 4344
rect 1765 4340 1769 4344
rect 1785 4340 1789 4344
rect 1831 4340 1835 4344
rect 1905 4340 1909 4344
rect 1951 4340 1955 4344
rect 1971 4340 1975 4344
rect 1991 4340 1995 4344
rect 2051 4340 2055 4344
rect 2059 4340 2063 4344
rect 2131 4340 2135 4344
rect 2196 4340 2200 4344
rect 2204 4340 2208 4344
rect 2226 4340 2230 4344
rect 2315 4340 2319 4344
rect 2325 4340 2329 4344
rect 2355 4340 2359 4344
rect 2365 4340 2369 4344
rect 2411 4340 2415 4344
rect 2421 4340 2425 4344
rect 2441 4340 2445 4344
rect 2511 4340 2515 4344
rect 2531 4340 2535 4344
rect 2551 4340 2555 4344
rect 2625 4340 2629 4344
rect 2645 4340 2649 4344
rect 2665 4340 2669 4344
rect 2685 4340 2689 4344
rect 2735 4340 2739 4344
rect 2755 4340 2759 4344
rect 2769 4340 2773 4344
rect 2789 4340 2793 4344
rect 2801 4340 2805 4344
rect 2821 4340 2825 4344
rect 2867 4340 2871 4344
rect 2875 4340 2879 4344
rect 2895 4340 2899 4344
rect 2903 4340 2907 4344
rect 2925 4340 2929 4344
rect 2985 4340 2989 4344
rect 3050 4340 3054 4344
rect 3072 4340 3076 4344
rect 3080 4340 3084 4344
rect 3157 4340 3161 4344
rect 3165 4340 3169 4344
rect 3230 4340 3234 4344
rect 3252 4340 3256 4344
rect 3260 4340 3264 4344
rect 3337 4340 3341 4344
rect 3345 4340 3349 4344
rect 3405 4340 3409 4344
rect 3451 4340 3455 4344
rect 3473 4340 3477 4344
rect 3481 4340 3485 4344
rect 3501 4340 3505 4344
rect 3509 4340 3513 4344
rect 3555 4340 3559 4344
rect 3575 4340 3579 4344
rect 3587 4340 3591 4344
rect 3607 4340 3611 4344
rect 3621 4340 3625 4344
rect 3641 4340 3645 4344
rect 3696 4340 3700 4344
rect 3704 4340 3708 4344
rect 3726 4340 3730 4344
rect 3791 4340 3795 4344
rect 3811 4340 3815 4344
rect 3885 4340 3889 4344
rect 3905 4340 3909 4344
rect 3925 4340 3929 4344
rect 3945 4340 3949 4344
rect 3965 4340 3969 4344
rect 3985 4340 3989 4344
rect 4005 4340 4009 4344
rect 4025 4340 4029 4344
rect 4083 4340 4087 4344
rect 4105 4340 4109 4344
rect 4151 4340 4155 4344
rect 4171 4340 4175 4344
rect 4231 4340 4235 4344
rect 4296 4340 4300 4344
rect 4304 4340 4308 4344
rect 4326 4340 4330 4344
rect 4391 4340 4395 4344
rect 4413 4340 4417 4344
rect 4421 4340 4425 4344
rect 4441 4340 4445 4344
rect 4449 4340 4453 4344
rect 4495 4340 4499 4344
rect 4515 4340 4519 4344
rect 4527 4340 4531 4344
rect 4547 4340 4551 4344
rect 4561 4340 4565 4344
rect 4581 4340 4585 4344
rect 4631 4340 4635 4344
rect 4653 4340 4657 4344
rect 4711 4340 4715 4344
rect 4731 4340 4735 4344
rect 45 4316 49 4320
rect 65 4316 69 4320
rect 111 4316 115 4320
rect 131 4316 135 4320
rect 151 4316 155 4320
rect 225 4316 229 4320
rect 245 4316 249 4320
rect 317 4316 321 4320
rect 325 4316 329 4320
rect 390 4316 394 4320
rect 412 4316 416 4320
rect 420 4316 424 4320
rect 476 4316 480 4320
rect 484 4316 488 4320
rect 506 4316 510 4320
rect 585 4316 589 4320
rect 645 4316 649 4320
rect 665 4316 669 4320
rect 685 4316 689 4320
rect 745 4316 749 4320
rect 791 4316 795 4320
rect 811 4316 815 4320
rect 831 4316 835 4320
rect 905 4316 909 4320
rect 925 4316 929 4320
rect 945 4316 949 4320
rect 965 4316 969 4320
rect 1025 4316 1029 4320
rect 1045 4316 1049 4320
rect 1065 4316 1069 4320
rect 1111 4316 1115 4320
rect 1131 4316 1135 4320
rect 1151 4316 1155 4320
rect 1225 4316 1229 4320
rect 1245 4316 1249 4320
rect 1305 4316 1309 4320
rect 1325 4316 1329 4320
rect 1345 4316 1349 4320
rect 1405 4316 1409 4320
rect 1425 4316 1429 4320
rect 1471 4316 1475 4320
rect 1491 4316 1495 4320
rect 1511 4316 1515 4320
rect 1597 4316 1601 4320
rect 1605 4316 1609 4320
rect 1677 4316 1681 4320
rect 1685 4316 1689 4320
rect 1736 4316 1740 4320
rect 1744 4316 1748 4320
rect 1766 4316 1770 4320
rect 1845 4316 1849 4320
rect 1865 4316 1869 4320
rect 1911 4316 1915 4320
rect 1971 4316 1975 4320
rect 1991 4316 1995 4320
rect 2011 4316 2015 4320
rect 2071 4316 2075 4320
rect 2091 4316 2095 4320
rect 2111 4316 2115 4320
rect 2175 4316 2179 4320
rect 2195 4316 2199 4320
rect 2209 4316 2213 4320
rect 2229 4316 2233 4320
rect 2241 4316 2245 4320
rect 2261 4316 2265 4320
rect 2307 4316 2311 4320
rect 2315 4316 2319 4320
rect 2335 4316 2339 4320
rect 2343 4316 2347 4320
rect 2365 4316 2369 4320
rect 2411 4316 2415 4320
rect 2433 4316 2437 4320
rect 2505 4316 2509 4320
rect 2577 4316 2581 4320
rect 2585 4316 2589 4320
rect 2631 4316 2635 4320
rect 2653 4316 2657 4320
rect 2661 4316 2665 4320
rect 2681 4316 2685 4320
rect 2689 4316 2693 4320
rect 2735 4316 2739 4320
rect 2755 4316 2759 4320
rect 2767 4316 2771 4320
rect 2787 4316 2791 4320
rect 2801 4316 2805 4320
rect 2821 4316 2825 4320
rect 2871 4316 2875 4320
rect 2957 4316 2961 4320
rect 2965 4316 2969 4320
rect 3016 4316 3020 4320
rect 3024 4316 3028 4320
rect 3046 4316 3050 4320
rect 3111 4316 3115 4320
rect 3131 4316 3135 4320
rect 3205 4316 3209 4320
rect 3225 4316 3229 4320
rect 3285 4316 3289 4320
rect 3305 4316 3309 4320
rect 3351 4316 3355 4320
rect 3359 4316 3363 4320
rect 3435 4316 3439 4320
rect 3455 4316 3459 4320
rect 3469 4316 3473 4320
rect 3489 4316 3493 4320
rect 3501 4316 3505 4320
rect 3521 4316 3525 4320
rect 3567 4316 3571 4320
rect 3575 4316 3579 4320
rect 3595 4316 3599 4320
rect 3603 4316 3607 4320
rect 3625 4316 3629 4320
rect 3685 4316 3689 4320
rect 3705 4316 3709 4320
rect 3751 4316 3755 4320
rect 3759 4316 3763 4320
rect 3831 4316 3835 4320
rect 3853 4316 3857 4320
rect 3861 4316 3865 4320
rect 3881 4316 3885 4320
rect 3889 4316 3893 4320
rect 3935 4316 3939 4320
rect 3955 4316 3959 4320
rect 3967 4316 3971 4320
rect 3987 4316 3991 4320
rect 4001 4316 4005 4320
rect 4021 4316 4025 4320
rect 4071 4316 4075 4320
rect 4079 4316 4083 4320
rect 4165 4316 4169 4320
rect 4185 4316 4189 4320
rect 4205 4316 4209 4320
rect 4251 4316 4255 4320
rect 4273 4316 4277 4320
rect 4357 4316 4361 4320
rect 4365 4316 4369 4320
rect 4425 4316 4429 4320
rect 4445 4316 4449 4320
rect 4465 4316 4469 4320
rect 4511 4316 4515 4320
rect 4533 4316 4537 4320
rect 4541 4316 4545 4320
rect 4561 4316 4565 4320
rect 4569 4316 4573 4320
rect 4615 4316 4619 4320
rect 4635 4316 4639 4320
rect 4647 4316 4651 4320
rect 4667 4316 4671 4320
rect 4681 4316 4685 4320
rect 4701 4316 4705 4320
rect 45 4199 49 4276
rect 46 4187 49 4199
rect 43 4171 49 4187
rect 65 4199 69 4276
rect 111 4222 115 4236
rect 131 4222 135 4236
rect 99 4216 115 4222
rect 120 4216 135 4222
rect 65 4187 74 4199
rect 65 4171 71 4187
rect 99 4179 106 4216
rect 120 4193 126 4216
rect 43 4164 57 4171
rect 53 4144 57 4164
rect 63 4164 71 4171
rect 63 4144 67 4164
rect 99 4154 106 4167
rect 99 4148 118 4154
rect 114 4144 118 4148
rect 122 4144 126 4181
rect 151 4179 155 4236
rect 225 4199 229 4276
rect 226 4187 229 4199
rect 146 4167 155 4179
rect 223 4171 229 4187
rect 245 4199 249 4276
rect 317 4213 321 4236
rect 306 4201 321 4213
rect 325 4213 329 4236
rect 390 4233 394 4276
rect 387 4221 394 4233
rect 325 4201 334 4213
rect 245 4187 254 4199
rect 245 4171 251 4187
rect 144 4124 148 4167
rect 223 4164 237 4171
rect 233 4144 237 4164
rect 243 4164 251 4171
rect 243 4144 247 4164
rect 305 4124 309 4201
rect 325 4124 329 4201
rect 385 4144 389 4221
rect 412 4179 416 4236
rect 420 4232 424 4236
rect 476 4232 480 4236
rect 420 4224 438 4232
rect 434 4213 438 4224
rect 462 4224 480 4232
rect 462 4213 466 4224
rect 405 4167 414 4179
rect 405 4144 409 4167
rect 434 4156 438 4201
rect 425 4149 438 4156
rect 462 4156 466 4201
rect 484 4179 488 4236
rect 506 4233 510 4276
rect 506 4221 513 4233
rect 486 4167 495 4179
rect 462 4149 475 4156
rect 425 4144 429 4149
rect 471 4144 475 4149
rect 491 4144 495 4167
rect 511 4144 515 4221
rect 585 4193 589 4276
rect 585 4181 594 4193
rect 585 4124 589 4181
rect 645 4179 649 4236
rect 665 4222 669 4236
rect 685 4222 689 4236
rect 665 4216 680 4222
rect 685 4216 701 4222
rect 674 4193 680 4216
rect 645 4167 654 4179
rect 652 4124 656 4167
rect 674 4144 678 4181
rect 694 4179 701 4216
rect 745 4193 749 4276
rect 791 4268 795 4276
rect 780 4264 795 4268
rect 811 4264 815 4276
rect 780 4233 786 4264
rect 800 4260 815 4264
rect 800 4253 806 4260
rect 786 4221 796 4233
rect 745 4181 754 4193
rect 694 4154 701 4167
rect 682 4148 701 4154
rect 682 4144 686 4148
rect 745 4124 749 4181
rect 792 4164 796 4221
rect 800 4164 804 4241
rect 831 4233 835 4276
rect 808 4221 815 4233
rect 827 4221 835 4233
rect 808 4164 812 4221
rect 905 4213 909 4236
rect 906 4201 909 4213
rect 900 4153 906 4201
rect 925 4179 929 4236
rect 945 4214 949 4236
rect 965 4214 969 4236
rect 1025 4233 1029 4276
rect 1045 4264 1049 4276
rect 1065 4268 1069 4276
rect 1111 4268 1115 4276
rect 1065 4264 1080 4268
rect 1045 4260 1060 4264
rect 1054 4253 1060 4260
rect 1025 4221 1033 4233
rect 1045 4221 1052 4233
rect 945 4208 958 4214
rect 965 4213 985 4214
rect 965 4208 973 4213
rect 954 4179 958 4208
rect 927 4167 929 4179
rect 925 4165 929 4167
rect 925 4158 938 4165
rect 900 4149 930 4153
rect 926 4144 930 4149
rect 934 4144 938 4158
rect 954 4144 958 4167
rect 973 4159 979 4201
rect 1048 4164 1052 4221
rect 1056 4164 1060 4241
rect 1074 4233 1080 4264
rect 1100 4264 1115 4268
rect 1131 4264 1135 4276
rect 1100 4233 1106 4264
rect 1120 4260 1135 4264
rect 1120 4253 1126 4260
rect 1064 4221 1074 4233
rect 1106 4221 1116 4233
rect 1064 4164 1068 4221
rect 1112 4164 1116 4221
rect 1120 4164 1124 4241
rect 1151 4233 1155 4276
rect 1128 4221 1135 4233
rect 1147 4221 1155 4233
rect 1128 4164 1132 4221
rect 1225 4199 1229 4276
rect 1226 4187 1229 4199
rect 1223 4171 1229 4187
rect 1245 4199 1249 4276
rect 1305 4233 1309 4276
rect 1325 4264 1329 4276
rect 1345 4268 1349 4276
rect 1345 4264 1360 4268
rect 1325 4260 1340 4264
rect 1334 4253 1340 4260
rect 1305 4221 1313 4233
rect 1325 4221 1332 4233
rect 1245 4187 1254 4199
rect 1245 4171 1251 4187
rect 1223 4164 1237 4171
rect 962 4152 979 4159
rect 962 4144 966 4152
rect 1233 4144 1237 4164
rect 1243 4164 1251 4171
rect 1328 4164 1332 4221
rect 1336 4164 1340 4241
rect 1354 4233 1360 4264
rect 1344 4221 1354 4233
rect 1344 4164 1348 4221
rect 1405 4199 1409 4276
rect 1406 4187 1409 4199
rect 1403 4171 1409 4187
rect 1425 4199 1429 4276
rect 1471 4268 1475 4276
rect 1460 4264 1475 4268
rect 1491 4264 1495 4276
rect 1460 4233 1466 4264
rect 1480 4260 1495 4264
rect 1480 4253 1486 4260
rect 1466 4221 1476 4233
rect 1425 4187 1434 4199
rect 1425 4171 1431 4187
rect 1403 4164 1417 4171
rect 1243 4144 1247 4164
rect 1413 4144 1417 4164
rect 1423 4164 1431 4171
rect 1472 4164 1476 4221
rect 1480 4164 1484 4241
rect 1511 4233 1515 4276
rect 1488 4221 1495 4233
rect 1507 4221 1515 4233
rect 1488 4164 1492 4221
rect 1597 4213 1601 4236
rect 1586 4201 1601 4213
rect 1605 4213 1609 4236
rect 1677 4213 1681 4236
rect 1605 4201 1614 4213
rect 1666 4201 1681 4213
rect 1685 4213 1689 4236
rect 1736 4232 1740 4236
rect 1722 4224 1740 4232
rect 1722 4213 1726 4224
rect 1685 4201 1694 4213
rect 1423 4144 1427 4164
rect 1585 4124 1589 4201
rect 1605 4124 1609 4201
rect 1665 4124 1669 4201
rect 1685 4124 1689 4201
rect 1722 4156 1726 4201
rect 1744 4179 1748 4236
rect 1766 4233 1770 4276
rect 1766 4221 1773 4233
rect 1746 4167 1755 4179
rect 1722 4149 1735 4156
rect 1731 4144 1735 4149
rect 1751 4144 1755 4167
rect 1771 4144 1775 4221
rect 1845 4199 1849 4276
rect 1846 4187 1849 4199
rect 1843 4171 1849 4187
rect 1865 4199 1869 4276
rect 1865 4187 1874 4199
rect 1911 4193 1915 4276
rect 1971 4268 1975 4276
rect 1960 4264 1975 4268
rect 1991 4264 1995 4276
rect 1960 4233 1966 4264
rect 1980 4260 1995 4264
rect 1980 4253 1986 4260
rect 1966 4221 1976 4233
rect 1865 4171 1871 4187
rect 1906 4181 1915 4193
rect 1843 4164 1857 4171
rect 1853 4144 1857 4164
rect 1863 4164 1871 4171
rect 1863 4144 1867 4164
rect 1911 4124 1915 4181
rect 1972 4164 1976 4221
rect 1980 4164 1984 4241
rect 2011 4233 2015 4276
rect 2071 4268 2075 4276
rect 2060 4264 2075 4268
rect 2091 4264 2095 4276
rect 2060 4233 2066 4264
rect 2080 4260 2095 4264
rect 2080 4253 2086 4260
rect 1988 4221 1995 4233
rect 2007 4221 2015 4233
rect 2066 4221 2076 4233
rect 1988 4164 1992 4221
rect 2072 4164 2076 4221
rect 2080 4164 2084 4241
rect 2111 4233 2115 4276
rect 2088 4221 2095 4233
rect 2107 4221 2115 4233
rect 2088 4164 2092 4221
rect 2175 4193 2179 4236
rect 2195 4194 2199 4276
rect 2209 4217 2213 4276
rect 2229 4236 2233 4276
rect 2241 4270 2245 4276
rect 2235 4224 2238 4236
rect 2209 4209 2218 4217
rect 2175 4144 2179 4181
rect 2195 4124 2199 4182
rect 2214 4180 2218 4209
rect 2234 4160 2238 4224
rect 2205 4156 2238 4160
rect 2205 4124 2209 4156
rect 2243 4148 2247 4258
rect 2261 4250 2265 4276
rect 2307 4272 2311 4276
rect 2275 4270 2311 4272
rect 2287 4268 2311 4270
rect 2229 4136 2231 4148
rect 2227 4124 2231 4136
rect 2237 4136 2239 4148
rect 2237 4124 2241 4136
rect 2259 4124 2263 4238
rect 2275 4132 2279 4258
rect 2315 4244 2319 4276
rect 2335 4256 2339 4296
rect 2343 4273 2347 4296
rect 2343 4266 2351 4273
rect 2313 4149 2319 4244
rect 2347 4237 2351 4266
rect 2343 4231 2351 4237
rect 2343 4185 2347 4231
rect 2365 4224 2369 4236
rect 2367 4212 2369 4224
rect 2411 4213 2415 4276
rect 2433 4230 2437 4236
rect 2435 4218 2437 4230
rect 2313 4145 2337 4149
rect 2299 4140 2317 4141
rect 2287 4136 2317 4140
rect 2275 4128 2309 4132
rect 2305 4124 2309 4128
rect 2313 4124 2317 4136
rect 2333 4124 2337 4145
rect 2343 4124 2347 4173
rect 2365 4144 2369 4212
rect 2406 4201 2415 4213
rect 2411 4124 2415 4201
rect 2505 4193 2509 4276
rect 2653 4273 2657 4296
rect 2649 4266 2657 4273
rect 2649 4237 2653 4266
rect 2661 4256 2665 4296
rect 2681 4244 2685 4276
rect 2689 4272 2693 4276
rect 2689 4270 2725 4272
rect 2689 4268 2713 4270
rect 2577 4213 2581 4236
rect 2566 4201 2581 4213
rect 2585 4213 2589 4236
rect 2631 4224 2635 4236
rect 2649 4231 2657 4237
rect 2585 4201 2594 4213
rect 2631 4212 2633 4224
rect 2505 4181 2514 4193
rect 2435 4150 2437 4162
rect 2433 4144 2437 4150
rect 2505 4124 2509 4181
rect 2565 4124 2569 4201
rect 2585 4124 2589 4201
rect 2631 4144 2635 4212
rect 2653 4185 2657 4231
rect 2653 4124 2657 4173
rect 2681 4149 2687 4244
rect 2663 4145 2687 4149
rect 2663 4124 2667 4145
rect 2683 4140 2701 4141
rect 2683 4136 2713 4140
rect 2683 4124 2687 4136
rect 2721 4132 2725 4258
rect 2735 4250 2739 4276
rect 2755 4270 2759 4276
rect 2691 4128 2725 4132
rect 2691 4124 2695 4128
rect 2737 4124 2741 4238
rect 2753 4148 2757 4258
rect 2767 4236 2771 4276
rect 2762 4224 2765 4236
rect 2762 4160 2766 4224
rect 2787 4217 2791 4276
rect 2782 4209 2791 4217
rect 2782 4180 2786 4209
rect 2801 4194 2805 4276
rect 2821 4193 2825 4236
rect 2871 4193 2875 4276
rect 2957 4213 2961 4236
rect 2946 4201 2961 4213
rect 2965 4213 2969 4236
rect 3016 4232 3020 4236
rect 3002 4224 3020 4232
rect 3002 4213 3006 4224
rect 2965 4201 2974 4213
rect 2762 4156 2795 4160
rect 2761 4136 2763 4148
rect 2759 4124 2763 4136
rect 2769 4136 2771 4148
rect 2769 4124 2773 4136
rect 2791 4124 2795 4156
rect 2801 4124 2805 4182
rect 2866 4181 2875 4193
rect 2821 4144 2825 4181
rect 2871 4124 2875 4181
rect 2945 4124 2949 4201
rect 2965 4124 2969 4201
rect 3002 4156 3006 4201
rect 3024 4179 3028 4236
rect 3046 4233 3050 4276
rect 3046 4221 3053 4233
rect 3026 4167 3035 4179
rect 3002 4149 3015 4156
rect 3011 4144 3015 4149
rect 3031 4144 3035 4167
rect 3051 4144 3055 4221
rect 3111 4199 3115 4276
rect 3106 4187 3115 4199
rect 3109 4171 3115 4187
rect 3131 4199 3135 4276
rect 3205 4199 3209 4276
rect 3131 4187 3134 4199
rect 3206 4187 3209 4199
rect 3131 4171 3137 4187
rect 3109 4164 3117 4171
rect 3113 4144 3117 4164
rect 3123 4164 3137 4171
rect 3203 4171 3209 4187
rect 3225 4199 3229 4276
rect 3285 4199 3289 4276
rect 3225 4187 3234 4199
rect 3286 4187 3289 4199
rect 3225 4171 3231 4187
rect 3203 4164 3217 4171
rect 3123 4144 3127 4164
rect 3213 4144 3217 4164
rect 3223 4164 3231 4171
rect 3283 4171 3289 4187
rect 3305 4199 3309 4276
rect 3351 4213 3355 4236
rect 3346 4201 3355 4213
rect 3359 4213 3363 4236
rect 3359 4201 3374 4213
rect 3305 4187 3314 4199
rect 3305 4171 3311 4187
rect 3283 4164 3297 4171
rect 3223 4144 3227 4164
rect 3293 4144 3297 4164
rect 3303 4164 3311 4171
rect 3303 4144 3307 4164
rect 3351 4124 3355 4201
rect 3371 4124 3375 4201
rect 3435 4193 3439 4236
rect 3455 4194 3459 4276
rect 3469 4217 3473 4276
rect 3489 4236 3493 4276
rect 3501 4270 3505 4276
rect 3495 4224 3498 4236
rect 3469 4209 3478 4217
rect 3435 4144 3439 4181
rect 3455 4124 3459 4182
rect 3474 4180 3478 4209
rect 3494 4160 3498 4224
rect 3465 4156 3498 4160
rect 3465 4124 3469 4156
rect 3503 4148 3507 4258
rect 3521 4250 3525 4276
rect 3567 4272 3571 4276
rect 3535 4270 3571 4272
rect 3547 4268 3571 4270
rect 3489 4136 3491 4148
rect 3487 4124 3491 4136
rect 3497 4136 3499 4148
rect 3497 4124 3501 4136
rect 3519 4124 3523 4238
rect 3535 4132 3539 4258
rect 3575 4244 3579 4276
rect 3595 4256 3599 4296
rect 3603 4273 3607 4296
rect 3603 4266 3611 4273
rect 3573 4149 3579 4244
rect 3607 4237 3611 4266
rect 3603 4231 3611 4237
rect 3603 4185 3607 4231
rect 3625 4224 3629 4236
rect 3627 4212 3629 4224
rect 3573 4145 3597 4149
rect 3559 4140 3577 4141
rect 3547 4136 3577 4140
rect 3535 4128 3569 4132
rect 3565 4124 3569 4128
rect 3573 4124 3577 4136
rect 3593 4124 3597 4145
rect 3603 4124 3607 4173
rect 3625 4144 3629 4212
rect 3685 4199 3689 4276
rect 3686 4187 3689 4199
rect 3683 4171 3689 4187
rect 3705 4199 3709 4276
rect 3853 4273 3857 4296
rect 3849 4266 3857 4273
rect 3849 4237 3853 4266
rect 3861 4256 3865 4296
rect 3881 4244 3885 4276
rect 3889 4272 3893 4276
rect 3889 4270 3925 4272
rect 3889 4268 3913 4270
rect 3751 4213 3755 4236
rect 3746 4201 3755 4213
rect 3759 4213 3763 4236
rect 3831 4224 3835 4236
rect 3849 4231 3857 4237
rect 3759 4201 3774 4213
rect 3831 4212 3833 4224
rect 3705 4187 3714 4199
rect 3705 4171 3711 4187
rect 3683 4164 3697 4171
rect 3693 4144 3697 4164
rect 3703 4164 3711 4171
rect 3703 4144 3707 4164
rect 3751 4124 3755 4201
rect 3771 4124 3775 4201
rect 3831 4144 3835 4212
rect 3853 4185 3857 4231
rect 3853 4124 3857 4173
rect 3881 4149 3887 4244
rect 3863 4145 3887 4149
rect 3863 4124 3867 4145
rect 3883 4140 3901 4141
rect 3883 4136 3913 4140
rect 3883 4124 3887 4136
rect 3921 4132 3925 4258
rect 3935 4250 3939 4276
rect 3955 4270 3959 4276
rect 3891 4128 3925 4132
rect 3891 4124 3895 4128
rect 3937 4124 3941 4238
rect 3953 4148 3957 4258
rect 3967 4236 3971 4276
rect 3962 4224 3965 4236
rect 3962 4160 3966 4224
rect 3987 4217 3991 4276
rect 3982 4209 3991 4217
rect 3982 4180 3986 4209
rect 4001 4194 4005 4276
rect 4021 4193 4025 4236
rect 4071 4213 4075 4236
rect 4066 4201 4075 4213
rect 4079 4213 4083 4236
rect 4079 4201 4094 4213
rect 3962 4156 3995 4160
rect 3961 4136 3963 4148
rect 3959 4124 3963 4136
rect 3969 4136 3971 4148
rect 3969 4124 3973 4136
rect 3991 4124 3995 4156
rect 4001 4124 4005 4182
rect 4021 4144 4025 4181
rect 4071 4124 4075 4201
rect 4091 4124 4095 4201
rect 4165 4179 4169 4236
rect 4185 4222 4189 4236
rect 4205 4222 4209 4236
rect 4185 4216 4200 4222
rect 4205 4216 4221 4222
rect 4194 4193 4200 4216
rect 4165 4167 4174 4179
rect 4172 4124 4176 4167
rect 4194 4144 4198 4181
rect 4214 4179 4221 4216
rect 4251 4213 4255 4276
rect 4533 4273 4537 4296
rect 4529 4266 4537 4273
rect 4529 4237 4533 4266
rect 4541 4256 4545 4296
rect 4561 4244 4565 4276
rect 4569 4272 4573 4276
rect 4569 4270 4605 4272
rect 4569 4268 4593 4270
rect 4273 4230 4277 4236
rect 4275 4218 4277 4230
rect 4357 4213 4361 4236
rect 4246 4201 4255 4213
rect 4346 4201 4361 4213
rect 4365 4213 4369 4236
rect 4365 4201 4374 4213
rect 4214 4154 4221 4167
rect 4202 4148 4221 4154
rect 4202 4144 4206 4148
rect 4251 4124 4255 4201
rect 4275 4150 4277 4162
rect 4273 4144 4277 4150
rect 4345 4124 4349 4201
rect 4365 4124 4369 4201
rect 4425 4179 4429 4236
rect 4445 4222 4449 4236
rect 4465 4222 4469 4236
rect 4511 4224 4515 4236
rect 4529 4231 4537 4237
rect 4445 4216 4460 4222
rect 4465 4216 4481 4222
rect 4454 4193 4460 4216
rect 4425 4167 4434 4179
rect 4432 4124 4436 4167
rect 4454 4144 4458 4181
rect 4474 4179 4481 4216
rect 4511 4212 4513 4224
rect 4474 4154 4481 4167
rect 4462 4148 4481 4154
rect 4462 4144 4466 4148
rect 4511 4144 4515 4212
rect 4533 4185 4537 4231
rect 4533 4124 4537 4173
rect 4561 4149 4567 4244
rect 4543 4145 4567 4149
rect 4543 4124 4547 4145
rect 4563 4140 4581 4141
rect 4563 4136 4593 4140
rect 4563 4124 4567 4136
rect 4601 4132 4605 4258
rect 4615 4250 4619 4276
rect 4635 4270 4639 4276
rect 4571 4128 4605 4132
rect 4571 4124 4575 4128
rect 4617 4124 4621 4238
rect 4633 4148 4637 4258
rect 4647 4236 4651 4276
rect 4642 4224 4645 4236
rect 4642 4160 4646 4224
rect 4667 4217 4671 4276
rect 4662 4209 4671 4217
rect 4662 4180 4666 4209
rect 4681 4194 4685 4276
rect 4701 4193 4705 4236
rect 4642 4156 4675 4160
rect 4641 4136 4643 4148
rect 4639 4124 4643 4136
rect 4649 4136 4651 4148
rect 4649 4124 4653 4136
rect 4671 4124 4675 4156
rect 4681 4124 4685 4182
rect 4701 4144 4705 4181
rect 53 4100 57 4104
rect 63 4100 67 4104
rect 114 4100 118 4104
rect 122 4100 126 4104
rect 144 4100 148 4104
rect 233 4100 237 4104
rect 243 4100 247 4104
rect 305 4100 309 4104
rect 325 4100 329 4104
rect 385 4100 389 4104
rect 405 4100 409 4104
rect 425 4100 429 4104
rect 471 4100 475 4104
rect 491 4100 495 4104
rect 511 4100 515 4104
rect 585 4100 589 4104
rect 652 4100 656 4104
rect 674 4100 678 4104
rect 682 4100 686 4104
rect 745 4100 749 4104
rect 792 4100 796 4104
rect 800 4100 804 4104
rect 808 4100 812 4104
rect 926 4100 930 4104
rect 934 4100 938 4104
rect 954 4100 958 4104
rect 962 4100 966 4104
rect 1048 4100 1052 4104
rect 1056 4100 1060 4104
rect 1064 4100 1068 4104
rect 1112 4100 1116 4104
rect 1120 4100 1124 4104
rect 1128 4100 1132 4104
rect 1233 4100 1237 4104
rect 1243 4100 1247 4104
rect 1328 4100 1332 4104
rect 1336 4100 1340 4104
rect 1344 4100 1348 4104
rect 1413 4100 1417 4104
rect 1423 4100 1427 4104
rect 1472 4100 1476 4104
rect 1480 4100 1484 4104
rect 1488 4100 1492 4104
rect 1585 4100 1589 4104
rect 1605 4100 1609 4104
rect 1665 4100 1669 4104
rect 1685 4100 1689 4104
rect 1731 4100 1735 4104
rect 1751 4100 1755 4104
rect 1771 4100 1775 4104
rect 1853 4100 1857 4104
rect 1863 4100 1867 4104
rect 1911 4100 1915 4104
rect 1972 4100 1976 4104
rect 1980 4100 1984 4104
rect 1988 4100 1992 4104
rect 2072 4100 2076 4104
rect 2080 4100 2084 4104
rect 2088 4100 2092 4104
rect 2175 4100 2179 4104
rect 2195 4100 2199 4104
rect 2205 4100 2209 4104
rect 2227 4100 2231 4104
rect 2237 4100 2241 4104
rect 2259 4100 2263 4104
rect 2305 4100 2309 4104
rect 2313 4100 2317 4104
rect 2333 4100 2337 4104
rect 2343 4100 2347 4104
rect 2365 4100 2369 4104
rect 2411 4100 2415 4104
rect 2433 4100 2437 4104
rect 2505 4100 2509 4104
rect 2565 4100 2569 4104
rect 2585 4100 2589 4104
rect 2631 4100 2635 4104
rect 2653 4100 2657 4104
rect 2663 4100 2667 4104
rect 2683 4100 2687 4104
rect 2691 4100 2695 4104
rect 2737 4100 2741 4104
rect 2759 4100 2763 4104
rect 2769 4100 2773 4104
rect 2791 4100 2795 4104
rect 2801 4100 2805 4104
rect 2821 4100 2825 4104
rect 2871 4100 2875 4104
rect 2945 4100 2949 4104
rect 2965 4100 2969 4104
rect 3011 4100 3015 4104
rect 3031 4100 3035 4104
rect 3051 4100 3055 4104
rect 3113 4100 3117 4104
rect 3123 4100 3127 4104
rect 3213 4100 3217 4104
rect 3223 4100 3227 4104
rect 3293 4100 3297 4104
rect 3303 4100 3307 4104
rect 3351 4100 3355 4104
rect 3371 4100 3375 4104
rect 3435 4100 3439 4104
rect 3455 4100 3459 4104
rect 3465 4100 3469 4104
rect 3487 4100 3491 4104
rect 3497 4100 3501 4104
rect 3519 4100 3523 4104
rect 3565 4100 3569 4104
rect 3573 4100 3577 4104
rect 3593 4100 3597 4104
rect 3603 4100 3607 4104
rect 3625 4100 3629 4104
rect 3693 4100 3697 4104
rect 3703 4100 3707 4104
rect 3751 4100 3755 4104
rect 3771 4100 3775 4104
rect 3831 4100 3835 4104
rect 3853 4100 3857 4104
rect 3863 4100 3867 4104
rect 3883 4100 3887 4104
rect 3891 4100 3895 4104
rect 3937 4100 3941 4104
rect 3959 4100 3963 4104
rect 3969 4100 3973 4104
rect 3991 4100 3995 4104
rect 4001 4100 4005 4104
rect 4021 4100 4025 4104
rect 4071 4100 4075 4104
rect 4091 4100 4095 4104
rect 4172 4100 4176 4104
rect 4194 4100 4198 4104
rect 4202 4100 4206 4104
rect 4251 4100 4255 4104
rect 4273 4100 4277 4104
rect 4345 4100 4349 4104
rect 4365 4100 4369 4104
rect 4432 4100 4436 4104
rect 4454 4100 4458 4104
rect 4462 4100 4466 4104
rect 4511 4100 4515 4104
rect 4533 4100 4537 4104
rect 4543 4100 4547 4104
rect 4563 4100 4567 4104
rect 4571 4100 4575 4104
rect 4617 4100 4621 4104
rect 4639 4100 4643 4104
rect 4649 4100 4653 4104
rect 4671 4100 4675 4104
rect 4681 4100 4685 4104
rect 4701 4100 4705 4104
rect 53 4076 57 4080
rect 63 4076 67 4080
rect 113 4076 117 4080
rect 123 4076 127 4080
rect 213 4076 217 4080
rect 223 4076 227 4080
rect 285 4076 289 4080
rect 305 4076 309 4080
rect 325 4076 329 4080
rect 374 4076 378 4080
rect 382 4076 386 4080
rect 404 4076 408 4080
rect 485 4076 489 4080
rect 505 4076 509 4080
rect 553 4076 557 4080
rect 563 4076 567 4080
rect 631 4076 635 4080
rect 651 4076 655 4080
rect 671 4076 675 4080
rect 768 4076 772 4080
rect 776 4076 780 4080
rect 784 4076 788 4080
rect 832 4076 836 4080
rect 840 4076 844 4080
rect 848 4076 852 4080
rect 945 4076 949 4080
rect 965 4076 969 4080
rect 985 4076 989 4080
rect 1031 4076 1035 4080
rect 1051 4076 1055 4080
rect 1071 4076 1075 4080
rect 1145 4076 1149 4080
rect 1228 4076 1232 4080
rect 1236 4076 1240 4080
rect 1244 4076 1248 4080
rect 1291 4076 1295 4080
rect 1352 4076 1356 4080
rect 1360 4076 1364 4080
rect 1368 4076 1372 4080
rect 1452 4076 1456 4080
rect 1460 4076 1464 4080
rect 1468 4076 1472 4080
rect 1553 4076 1557 4080
rect 1563 4076 1567 4080
rect 1645 4076 1649 4080
rect 1665 4076 1669 4080
rect 1735 4076 1739 4080
rect 1755 4076 1759 4080
rect 1765 4076 1769 4080
rect 1825 4076 1829 4080
rect 1845 4076 1849 4080
rect 1865 4076 1869 4080
rect 1911 4076 1915 4080
rect 1931 4076 1935 4080
rect 2005 4076 2009 4080
rect 2051 4076 2055 4080
rect 2071 4076 2075 4080
rect 2091 4076 2095 4080
rect 2151 4076 2155 4080
rect 2213 4076 2217 4080
rect 2223 4076 2227 4080
rect 2292 4076 2296 4080
rect 2300 4076 2304 4080
rect 2308 4076 2312 4080
rect 2391 4076 2395 4080
rect 2413 4076 2417 4080
rect 2471 4076 2475 4080
rect 2491 4076 2495 4080
rect 2511 4076 2515 4080
rect 2531 4076 2535 4080
rect 2551 4076 2555 4080
rect 2571 4076 2575 4080
rect 2591 4076 2595 4080
rect 2611 4076 2615 4080
rect 2675 4076 2679 4080
rect 2695 4076 2699 4080
rect 2705 4076 2709 4080
rect 2727 4076 2731 4080
rect 2737 4076 2741 4080
rect 2759 4076 2763 4080
rect 2805 4076 2809 4080
rect 2813 4076 2817 4080
rect 2833 4076 2837 4080
rect 2843 4076 2847 4080
rect 2865 4076 2869 4080
rect 2911 4076 2915 4080
rect 2971 4076 2975 4080
rect 2991 4076 2995 4080
rect 3011 4076 3015 4080
rect 3071 4076 3075 4080
rect 3091 4076 3095 4080
rect 3153 4076 3157 4080
rect 3163 4076 3167 4080
rect 3252 4076 3256 4080
rect 3274 4076 3278 4080
rect 3282 4076 3286 4080
rect 3331 4076 3335 4080
rect 3341 4076 3345 4080
rect 3361 4076 3365 4080
rect 3445 4076 3449 4080
rect 3465 4076 3469 4080
rect 3525 4076 3529 4080
rect 3571 4076 3575 4080
rect 3593 4076 3597 4080
rect 3603 4076 3607 4080
rect 3623 4076 3627 4080
rect 3631 4076 3635 4080
rect 3677 4076 3681 4080
rect 3699 4076 3703 4080
rect 3709 4076 3713 4080
rect 3731 4076 3735 4080
rect 3741 4076 3745 4080
rect 3761 4076 3765 4080
rect 3832 4076 3836 4080
rect 3854 4076 3858 4080
rect 3862 4076 3866 4080
rect 3911 4076 3915 4080
rect 3931 4076 3935 4080
rect 4005 4076 4009 4080
rect 4025 4076 4029 4080
rect 4071 4076 4075 4080
rect 4081 4076 4085 4080
rect 4101 4076 4105 4080
rect 4171 4076 4175 4080
rect 4191 4076 4195 4080
rect 4211 4076 4215 4080
rect 4285 4076 4289 4080
rect 4305 4076 4309 4080
rect 4325 4076 4329 4080
rect 4385 4076 4389 4080
rect 4431 4076 4435 4080
rect 4453 4076 4457 4080
rect 4463 4076 4467 4080
rect 4483 4076 4487 4080
rect 4491 4076 4495 4080
rect 4537 4076 4541 4080
rect 4559 4076 4563 4080
rect 4569 4076 4573 4080
rect 4591 4076 4595 4080
rect 4601 4076 4605 4080
rect 4621 4076 4625 4080
rect 4671 4076 4675 4080
rect 53 4016 57 4036
rect 43 4009 57 4016
rect 63 4016 67 4036
rect 113 4016 117 4036
rect 63 4009 71 4016
rect 43 3993 49 4009
rect 46 3981 49 3993
rect 45 3904 49 3981
rect 65 3993 71 4009
rect 109 4009 117 4016
rect 123 4016 127 4036
rect 213 4016 217 4036
rect 123 4009 137 4016
rect 109 3993 115 4009
rect 65 3981 74 3993
rect 106 3981 115 3993
rect 65 3904 69 3981
rect 111 3904 115 3981
rect 131 3993 137 4009
rect 203 4009 217 4016
rect 223 4016 227 4036
rect 223 4009 231 4016
rect 203 3993 209 4009
rect 131 3981 134 3993
rect 206 3981 209 3993
rect 131 3904 135 3981
rect 205 3904 209 3981
rect 225 3993 231 4009
rect 225 3981 234 3993
rect 225 3904 229 3981
rect 285 3959 289 4036
rect 305 4013 309 4036
rect 325 4031 329 4036
rect 374 4032 378 4036
rect 325 4024 338 4031
rect 305 4001 314 4013
rect 287 3947 294 3959
rect 290 3904 294 3947
rect 312 3944 316 4001
rect 334 3979 338 4024
rect 359 4026 378 4032
rect 359 4013 366 4026
rect 334 3956 338 3967
rect 359 3964 366 4001
rect 382 3999 386 4036
rect 404 4013 408 4056
rect 406 4001 415 4013
rect 380 3964 386 3987
rect 359 3958 375 3964
rect 380 3958 395 3964
rect 320 3948 338 3956
rect 320 3944 324 3948
rect 371 3944 375 3958
rect 391 3944 395 3958
rect 411 3944 415 4001
rect 485 3979 489 4056
rect 505 3979 509 4056
rect 553 4016 557 4036
rect 549 4009 557 4016
rect 563 4016 567 4036
rect 631 4031 635 4036
rect 622 4024 635 4031
rect 563 4009 577 4016
rect 549 3993 555 4009
rect 546 3981 555 3993
rect 486 3967 501 3979
rect 497 3944 501 3967
rect 505 3967 514 3979
rect 505 3944 509 3967
rect 551 3904 555 3981
rect 571 3993 577 4009
rect 571 3981 574 3993
rect 571 3904 575 3981
rect 622 3979 626 4024
rect 651 4013 655 4036
rect 646 4001 655 4013
rect 622 3956 626 3967
rect 622 3948 640 3956
rect 636 3944 640 3948
rect 644 3944 648 4001
rect 671 3959 675 4036
rect 768 3959 772 4016
rect 666 3947 673 3959
rect 745 3947 753 3959
rect 765 3947 772 3959
rect 666 3904 670 3947
rect 745 3904 749 3947
rect 776 3939 780 4016
rect 784 3959 788 4016
rect 832 3959 836 4016
rect 784 3947 794 3959
rect 826 3947 836 3959
rect 774 3920 780 3927
rect 765 3916 780 3920
rect 794 3916 800 3947
rect 765 3904 769 3916
rect 785 3912 800 3916
rect 820 3916 826 3947
rect 840 3939 844 4016
rect 848 3959 852 4016
rect 945 3959 949 4036
rect 965 4013 969 4036
rect 985 4031 989 4036
rect 1031 4031 1035 4036
rect 985 4024 998 4031
rect 965 4001 974 4013
rect 848 3947 855 3959
rect 867 3947 875 3959
rect 947 3947 954 3959
rect 840 3920 846 3927
rect 840 3916 855 3920
rect 820 3912 835 3916
rect 785 3904 789 3912
rect 831 3904 835 3912
rect 851 3904 855 3916
rect 871 3904 875 3947
rect 950 3904 954 3947
rect 972 3944 976 4001
rect 994 3979 998 4024
rect 1022 4024 1035 4031
rect 1022 3979 1026 4024
rect 1051 4013 1055 4036
rect 1046 4001 1055 4013
rect 994 3956 998 3967
rect 980 3948 998 3956
rect 1022 3956 1026 3967
rect 1022 3948 1040 3956
rect 980 3944 984 3948
rect 1036 3944 1040 3948
rect 1044 3944 1048 4001
rect 1071 3959 1075 4036
rect 1145 3999 1149 4056
rect 1145 3987 1154 3999
rect 1066 3947 1073 3959
rect 1066 3904 1070 3947
rect 1145 3904 1149 3987
rect 1228 3959 1232 4016
rect 1205 3947 1213 3959
rect 1225 3947 1232 3959
rect 1205 3904 1209 3947
rect 1236 3939 1240 4016
rect 1244 3959 1248 4016
rect 1291 3999 1295 4056
rect 1553 4016 1557 4036
rect 1286 3987 1295 3999
rect 1244 3947 1254 3959
rect 1234 3920 1240 3927
rect 1225 3916 1240 3920
rect 1254 3916 1260 3947
rect 1225 3904 1229 3916
rect 1245 3912 1260 3916
rect 1245 3904 1249 3912
rect 1291 3904 1295 3987
rect 1352 3959 1356 4016
rect 1346 3947 1356 3959
rect 1340 3916 1346 3947
rect 1360 3939 1364 4016
rect 1368 3959 1372 4016
rect 1452 3959 1456 4016
rect 1368 3947 1375 3959
rect 1387 3947 1395 3959
rect 1446 3947 1456 3959
rect 1360 3920 1366 3927
rect 1360 3916 1375 3920
rect 1340 3912 1355 3916
rect 1351 3904 1355 3912
rect 1371 3904 1375 3916
rect 1391 3904 1395 3947
rect 1440 3916 1446 3947
rect 1460 3939 1464 4016
rect 1468 3959 1472 4016
rect 1549 4009 1557 4016
rect 1563 4016 1567 4036
rect 1563 4009 1577 4016
rect 1549 3993 1555 4009
rect 1546 3981 1555 3993
rect 1468 3947 1475 3959
rect 1487 3947 1495 3959
rect 1460 3920 1466 3927
rect 1460 3916 1475 3920
rect 1440 3912 1455 3916
rect 1451 3904 1455 3912
rect 1471 3904 1475 3916
rect 1491 3904 1495 3947
rect 1551 3904 1555 3981
rect 1571 3993 1577 4009
rect 1571 3981 1574 3993
rect 1571 3904 1575 3981
rect 1645 3979 1649 4056
rect 1665 3979 1669 4056
rect 1735 4030 1739 4036
rect 1721 4018 1733 4030
rect 1646 3967 1661 3979
rect 1657 3944 1661 3967
rect 1665 3967 1674 3979
rect 1665 3944 1669 3967
rect 1721 3944 1725 4018
rect 1755 3993 1759 4036
rect 1746 3981 1759 3993
rect 1743 3904 1747 3981
rect 1765 3979 1769 4036
rect 1765 3967 1774 3979
rect 1765 3904 1769 3967
rect 1825 3959 1829 4036
rect 1845 4013 1849 4036
rect 1865 4031 1869 4036
rect 1865 4024 1878 4031
rect 1845 4001 1854 4013
rect 1827 3947 1834 3959
rect 1830 3904 1834 3947
rect 1852 3944 1856 4001
rect 1874 3979 1878 4024
rect 1911 3979 1915 4056
rect 1931 3979 1935 4056
rect 2005 3999 2009 4056
rect 2051 4031 2055 4036
rect 2042 4024 2055 4031
rect 2005 3987 2014 3999
rect 1906 3967 1915 3979
rect 1874 3956 1878 3967
rect 1860 3948 1878 3956
rect 1860 3944 1864 3948
rect 1911 3944 1915 3967
rect 1919 3967 1934 3979
rect 1919 3944 1923 3967
rect 2005 3904 2009 3987
rect 2042 3979 2046 4024
rect 2071 4013 2075 4036
rect 2066 4001 2075 4013
rect 2042 3956 2046 3967
rect 2042 3948 2060 3956
rect 2056 3944 2060 3948
rect 2064 3944 2068 4001
rect 2091 3959 2095 4036
rect 2151 3999 2155 4056
rect 2213 4016 2217 4036
rect 2146 3987 2155 3999
rect 2209 4009 2217 4016
rect 2223 4016 2227 4036
rect 2223 4009 2237 4016
rect 2209 3993 2215 4009
rect 2086 3947 2093 3959
rect 2086 3904 2090 3947
rect 2151 3904 2155 3987
rect 2206 3981 2215 3993
rect 2211 3904 2215 3981
rect 2231 3993 2237 4009
rect 2231 3981 2234 3993
rect 2231 3904 2235 3981
rect 2292 3959 2296 4016
rect 2286 3947 2296 3959
rect 2280 3916 2286 3947
rect 2300 3939 2304 4016
rect 2308 3959 2312 4016
rect 2391 3979 2395 4056
rect 2413 4030 2417 4036
rect 2415 4018 2417 4030
rect 2386 3967 2395 3979
rect 2308 3947 2315 3959
rect 2327 3947 2335 3959
rect 2300 3920 2306 3927
rect 2300 3916 2315 3920
rect 2280 3912 2295 3916
rect 2291 3904 2295 3912
rect 2311 3904 2315 3916
rect 2331 3904 2335 3947
rect 2391 3904 2395 3967
rect 2471 4013 2475 4036
rect 2491 4013 2495 4036
rect 2511 4016 2515 4036
rect 2531 4016 2535 4036
rect 2551 4016 2555 4036
rect 2571 4016 2575 4036
rect 2591 4016 2595 4036
rect 2611 4016 2615 4036
rect 2471 4001 2474 4013
rect 2486 4001 2495 4013
rect 2522 4004 2535 4016
rect 2562 4004 2575 4016
rect 2602 4004 2615 4016
rect 2415 3950 2417 3962
rect 2413 3944 2417 3950
rect 2471 3944 2475 4001
rect 2491 3944 2495 4001
rect 2511 3944 2515 4004
rect 2531 3944 2535 4004
rect 2551 3944 2555 4004
rect 2571 3944 2575 4004
rect 2591 3944 2595 4004
rect 2611 3944 2615 4004
rect 2675 3999 2679 4036
rect 2695 3998 2699 4056
rect 2705 4024 2709 4056
rect 2727 4044 2731 4056
rect 2729 4032 2731 4044
rect 2737 4044 2741 4056
rect 2737 4032 2739 4044
rect 2705 4020 2738 4024
rect 2675 3944 2679 3987
rect 2695 3904 2699 3986
rect 2714 3971 2718 4000
rect 2709 3963 2718 3971
rect 2709 3904 2713 3963
rect 2734 3956 2738 4020
rect 2735 3944 2738 3956
rect 2729 3904 2733 3944
rect 2743 3922 2747 4032
rect 2759 3942 2763 4056
rect 2805 4052 2809 4056
rect 2775 4048 2809 4052
rect 2741 3904 2745 3910
rect 2761 3904 2765 3930
rect 2775 3922 2779 4048
rect 2813 4044 2817 4056
rect 2787 4040 2817 4044
rect 2799 4039 2817 4040
rect 2833 4035 2837 4056
rect 2813 4031 2837 4035
rect 2813 3936 2819 4031
rect 2843 4007 2847 4056
rect 2843 3949 2847 3995
rect 2865 3968 2869 4036
rect 2911 3999 2915 4056
rect 2971 4031 2975 4036
rect 2906 3987 2915 3999
rect 2867 3956 2869 3968
rect 2843 3943 2851 3949
rect 2865 3944 2869 3956
rect 2787 3910 2811 3912
rect 2775 3908 2811 3910
rect 2807 3904 2811 3908
rect 2815 3904 2819 3936
rect 2835 3884 2839 3924
rect 2847 3914 2851 3943
rect 2843 3907 2851 3914
rect 2843 3884 2847 3907
rect 2911 3904 2915 3987
rect 2962 4024 2975 4031
rect 2962 3979 2966 4024
rect 2991 4013 2995 4036
rect 2986 4001 2995 4013
rect 2962 3956 2966 3967
rect 2962 3948 2980 3956
rect 2976 3944 2980 3948
rect 2984 3944 2988 4001
rect 3011 3959 3015 4036
rect 3071 3979 3075 4056
rect 3091 3979 3095 4056
rect 3153 4016 3157 4036
rect 3149 4009 3157 4016
rect 3163 4016 3167 4036
rect 3163 4009 3177 4016
rect 3252 4013 3256 4056
rect 3149 3993 3155 4009
rect 3146 3981 3155 3993
rect 3066 3967 3075 3979
rect 3006 3947 3013 3959
rect 3006 3904 3010 3947
rect 3071 3944 3075 3967
rect 3079 3967 3094 3979
rect 3079 3944 3083 3967
rect 3151 3904 3155 3981
rect 3171 3993 3177 4009
rect 3245 4001 3254 4013
rect 3171 3981 3174 3993
rect 3171 3904 3175 3981
rect 3245 3944 3249 4001
rect 3274 3999 3278 4036
rect 3282 4032 3286 4036
rect 3282 4026 3301 4032
rect 3294 4013 3301 4026
rect 3274 3964 3280 3987
rect 3294 3964 3301 4001
rect 3331 3979 3335 4036
rect 3341 3993 3345 4036
rect 3361 4030 3365 4036
rect 3367 4018 3379 4030
rect 3341 3981 3354 3993
rect 3326 3967 3335 3979
rect 3265 3958 3280 3964
rect 3285 3958 3301 3964
rect 3265 3944 3269 3958
rect 3285 3944 3289 3958
rect 3331 3904 3335 3967
rect 3353 3904 3357 3981
rect 3375 3944 3379 4018
rect 3445 3979 3449 4056
rect 3465 3979 3469 4056
rect 3525 3999 3529 4056
rect 3525 3987 3534 3999
rect 3446 3967 3461 3979
rect 3457 3944 3461 3967
rect 3465 3967 3474 3979
rect 3465 3944 3469 3967
rect 3525 3904 3529 3987
rect 3571 3968 3575 4036
rect 3593 4007 3597 4056
rect 3603 4035 3607 4056
rect 3623 4044 3627 4056
rect 3631 4052 3635 4056
rect 3631 4048 3665 4052
rect 3623 4040 3653 4044
rect 3623 4039 3641 4040
rect 3603 4031 3627 4035
rect 3571 3956 3573 3968
rect 3571 3944 3575 3956
rect 3593 3949 3597 3995
rect 3589 3943 3597 3949
rect 3589 3914 3593 3943
rect 3621 3936 3627 4031
rect 3589 3907 3597 3914
rect 3593 3884 3597 3907
rect 3601 3884 3605 3924
rect 3621 3904 3625 3936
rect 3661 3922 3665 4048
rect 3677 3942 3681 4056
rect 3699 4044 3703 4056
rect 3701 4032 3703 4044
rect 3709 4044 3713 4056
rect 3709 4032 3711 4044
rect 3629 3910 3653 3912
rect 3629 3908 3665 3910
rect 3629 3904 3633 3908
rect 3675 3904 3679 3930
rect 3693 3922 3697 4032
rect 3731 4024 3735 4056
rect 3702 4020 3735 4024
rect 3702 3956 3706 4020
rect 3722 3971 3726 4000
rect 3741 3998 3745 4056
rect 3761 3999 3765 4036
rect 3832 4013 3836 4056
rect 3825 4001 3834 4013
rect 3722 3963 3731 3971
rect 3702 3944 3705 3956
rect 3695 3904 3699 3910
rect 3707 3904 3711 3944
rect 3727 3904 3731 3963
rect 3741 3904 3745 3986
rect 3761 3944 3765 3987
rect 3825 3944 3829 4001
rect 3854 3999 3858 4036
rect 3862 4032 3866 4036
rect 3862 4026 3881 4032
rect 3874 4013 3881 4026
rect 3854 3964 3860 3987
rect 3874 3964 3881 4001
rect 3911 3979 3915 4056
rect 3931 3979 3935 4056
rect 4005 3979 4009 4056
rect 4025 3979 4029 4056
rect 4071 3979 4075 4036
rect 4081 3993 4085 4036
rect 4101 4030 4105 4036
rect 4171 4031 4175 4036
rect 4107 4018 4119 4030
rect 4081 3981 4094 3993
rect 3906 3967 3915 3979
rect 3845 3958 3860 3964
rect 3865 3958 3881 3964
rect 3845 3944 3849 3958
rect 3865 3944 3869 3958
rect 3911 3944 3915 3967
rect 3919 3967 3934 3979
rect 4006 3967 4021 3979
rect 3919 3944 3923 3967
rect 4017 3944 4021 3967
rect 4025 3967 4034 3979
rect 4066 3967 4075 3979
rect 4025 3944 4029 3967
rect 4071 3904 4075 3967
rect 4093 3904 4097 3981
rect 4115 3944 4119 4018
rect 4162 4024 4175 4031
rect 4162 3979 4166 4024
rect 4191 4013 4195 4036
rect 4186 4001 4195 4013
rect 4162 3956 4166 3967
rect 4162 3948 4180 3956
rect 4176 3944 4180 3948
rect 4184 3944 4188 4001
rect 4211 3959 4215 4036
rect 4285 3959 4289 4036
rect 4305 4013 4309 4036
rect 4325 4031 4329 4036
rect 4325 4024 4338 4031
rect 4305 4001 4314 4013
rect 4206 3947 4213 3959
rect 4287 3947 4294 3959
rect 4206 3904 4210 3947
rect 4290 3904 4294 3947
rect 4312 3944 4316 4001
rect 4334 3979 4338 4024
rect 4385 3999 4389 4056
rect 4385 3987 4394 3999
rect 4334 3956 4338 3967
rect 4320 3948 4338 3956
rect 4320 3944 4324 3948
rect 4385 3904 4389 3987
rect 4431 3968 4435 4036
rect 4453 4007 4457 4056
rect 4463 4035 4467 4056
rect 4483 4044 4487 4056
rect 4491 4052 4495 4056
rect 4491 4048 4525 4052
rect 4483 4040 4513 4044
rect 4483 4039 4501 4040
rect 4463 4031 4487 4035
rect 4431 3956 4433 3968
rect 4431 3944 4435 3956
rect 4453 3949 4457 3995
rect 4449 3943 4457 3949
rect 4449 3914 4453 3943
rect 4481 3936 4487 4031
rect 4449 3907 4457 3914
rect 4453 3884 4457 3907
rect 4461 3884 4465 3924
rect 4481 3904 4485 3936
rect 4521 3922 4525 4048
rect 4537 3942 4541 4056
rect 4559 4044 4563 4056
rect 4561 4032 4563 4044
rect 4569 4044 4573 4056
rect 4569 4032 4571 4044
rect 4489 3910 4513 3912
rect 4489 3908 4525 3910
rect 4489 3904 4493 3908
rect 4535 3904 4539 3930
rect 4553 3922 4557 4032
rect 4591 4024 4595 4056
rect 4562 4020 4595 4024
rect 4562 3956 4566 4020
rect 4582 3971 4586 4000
rect 4601 3998 4605 4056
rect 4621 3999 4625 4036
rect 4671 3999 4675 4056
rect 4666 3987 4675 3999
rect 4582 3963 4591 3971
rect 4562 3944 4565 3956
rect 4555 3904 4559 3910
rect 4567 3904 4571 3944
rect 4587 3904 4591 3963
rect 4601 3904 4605 3986
rect 4621 3944 4625 3987
rect 4671 3904 4675 3987
rect 45 3860 49 3864
rect 65 3860 69 3864
rect 111 3860 115 3864
rect 131 3860 135 3864
rect 205 3860 209 3864
rect 225 3860 229 3864
rect 290 3860 294 3864
rect 312 3860 316 3864
rect 320 3860 324 3864
rect 371 3860 375 3864
rect 391 3860 395 3864
rect 411 3860 415 3864
rect 497 3860 501 3864
rect 505 3860 509 3864
rect 551 3860 555 3864
rect 571 3860 575 3864
rect 636 3860 640 3864
rect 644 3860 648 3864
rect 666 3860 670 3864
rect 745 3860 749 3864
rect 765 3860 769 3864
rect 785 3860 789 3864
rect 831 3860 835 3864
rect 851 3860 855 3864
rect 871 3860 875 3864
rect 950 3860 954 3864
rect 972 3860 976 3864
rect 980 3860 984 3864
rect 1036 3860 1040 3864
rect 1044 3860 1048 3864
rect 1066 3860 1070 3864
rect 1145 3860 1149 3864
rect 1205 3860 1209 3864
rect 1225 3860 1229 3864
rect 1245 3860 1249 3864
rect 1291 3860 1295 3864
rect 1351 3860 1355 3864
rect 1371 3860 1375 3864
rect 1391 3860 1395 3864
rect 1451 3860 1455 3864
rect 1471 3860 1475 3864
rect 1491 3860 1495 3864
rect 1551 3860 1555 3864
rect 1571 3860 1575 3864
rect 1657 3860 1661 3864
rect 1665 3860 1669 3864
rect 1721 3860 1725 3864
rect 1743 3860 1747 3864
rect 1765 3860 1769 3864
rect 1830 3860 1834 3864
rect 1852 3860 1856 3864
rect 1860 3860 1864 3864
rect 1911 3860 1915 3864
rect 1919 3860 1923 3864
rect 2005 3860 2009 3864
rect 2056 3860 2060 3864
rect 2064 3860 2068 3864
rect 2086 3860 2090 3864
rect 2151 3860 2155 3864
rect 2211 3860 2215 3864
rect 2231 3860 2235 3864
rect 2291 3860 2295 3864
rect 2311 3860 2315 3864
rect 2331 3860 2335 3864
rect 2391 3860 2395 3864
rect 2413 3860 2417 3864
rect 2471 3860 2475 3864
rect 2491 3860 2495 3864
rect 2511 3860 2515 3864
rect 2531 3860 2535 3864
rect 2551 3860 2555 3864
rect 2571 3860 2575 3864
rect 2591 3860 2595 3864
rect 2611 3860 2615 3864
rect 2675 3860 2679 3864
rect 2695 3860 2699 3864
rect 2709 3860 2713 3864
rect 2729 3860 2733 3864
rect 2741 3860 2745 3864
rect 2761 3860 2765 3864
rect 2807 3860 2811 3864
rect 2815 3860 2819 3864
rect 2835 3860 2839 3864
rect 2843 3860 2847 3864
rect 2865 3860 2869 3864
rect 2911 3860 2915 3864
rect 2976 3860 2980 3864
rect 2984 3860 2988 3864
rect 3006 3860 3010 3864
rect 3071 3860 3075 3864
rect 3079 3860 3083 3864
rect 3151 3860 3155 3864
rect 3171 3860 3175 3864
rect 3245 3860 3249 3864
rect 3265 3860 3269 3864
rect 3285 3860 3289 3864
rect 3331 3860 3335 3864
rect 3353 3860 3357 3864
rect 3375 3860 3379 3864
rect 3457 3860 3461 3864
rect 3465 3860 3469 3864
rect 3525 3860 3529 3864
rect 3571 3860 3575 3864
rect 3593 3860 3597 3864
rect 3601 3860 3605 3864
rect 3621 3860 3625 3864
rect 3629 3860 3633 3864
rect 3675 3860 3679 3864
rect 3695 3860 3699 3864
rect 3707 3860 3711 3864
rect 3727 3860 3731 3864
rect 3741 3860 3745 3864
rect 3761 3860 3765 3864
rect 3825 3860 3829 3864
rect 3845 3860 3849 3864
rect 3865 3860 3869 3864
rect 3911 3860 3915 3864
rect 3919 3860 3923 3864
rect 4017 3860 4021 3864
rect 4025 3860 4029 3864
rect 4071 3860 4075 3864
rect 4093 3860 4097 3864
rect 4115 3860 4119 3864
rect 4176 3860 4180 3864
rect 4184 3860 4188 3864
rect 4206 3860 4210 3864
rect 4290 3860 4294 3864
rect 4312 3860 4316 3864
rect 4320 3860 4324 3864
rect 4385 3860 4389 3864
rect 4431 3860 4435 3864
rect 4453 3860 4457 3864
rect 4461 3860 4465 3864
rect 4481 3860 4485 3864
rect 4489 3860 4493 3864
rect 4535 3860 4539 3864
rect 4555 3860 4559 3864
rect 4567 3860 4571 3864
rect 4587 3860 4591 3864
rect 4601 3860 4605 3864
rect 4621 3860 4625 3864
rect 4671 3860 4675 3864
rect 57 3836 61 3840
rect 65 3836 69 3840
rect 116 3836 120 3840
rect 124 3836 128 3840
rect 146 3836 150 3840
rect 225 3836 229 3840
rect 285 3836 289 3840
rect 305 3836 309 3840
rect 325 3836 329 3840
rect 381 3836 385 3840
rect 403 3836 407 3840
rect 425 3836 429 3840
rect 485 3836 489 3840
rect 505 3836 509 3840
rect 565 3836 569 3840
rect 585 3836 589 3840
rect 631 3836 635 3840
rect 696 3836 700 3840
rect 704 3836 708 3840
rect 726 3836 730 3840
rect 791 3836 795 3840
rect 811 3836 815 3840
rect 885 3836 889 3840
rect 905 3836 909 3840
rect 925 3836 929 3840
rect 971 3836 975 3840
rect 991 3836 995 3840
rect 1011 3836 1015 3840
rect 1071 3836 1075 3840
rect 1091 3836 1095 3840
rect 1111 3836 1115 3840
rect 1171 3836 1175 3840
rect 1191 3836 1195 3840
rect 1211 3836 1215 3840
rect 1271 3836 1275 3840
rect 1345 3836 1349 3840
rect 1365 3836 1369 3840
rect 1385 3836 1389 3840
rect 1445 3836 1449 3840
rect 1510 3836 1514 3840
rect 1532 3836 1536 3840
rect 1540 3836 1544 3840
rect 1605 3836 1609 3840
rect 1651 3836 1655 3840
rect 1671 3836 1675 3840
rect 1691 3836 1695 3840
rect 1751 3836 1755 3840
rect 1759 3836 1763 3840
rect 1845 3836 1849 3840
rect 1865 3836 1869 3840
rect 1885 3836 1889 3840
rect 1945 3836 1949 3840
rect 1965 3836 1969 3840
rect 2011 3836 2015 3840
rect 2021 3836 2025 3840
rect 2041 3836 2045 3840
rect 2111 3836 2115 3840
rect 2133 3836 2137 3840
rect 2205 3836 2209 3840
rect 2225 3836 2229 3840
rect 2245 3836 2249 3840
rect 2265 3836 2269 3840
rect 2285 3836 2289 3840
rect 2305 3836 2309 3840
rect 2325 3836 2329 3840
rect 2345 3836 2349 3840
rect 2395 3836 2399 3840
rect 2415 3836 2419 3840
rect 2429 3836 2433 3840
rect 2449 3836 2453 3840
rect 2461 3836 2465 3840
rect 2481 3836 2485 3840
rect 2527 3836 2531 3840
rect 2535 3836 2539 3840
rect 2555 3836 2559 3840
rect 2563 3836 2567 3840
rect 2585 3836 2589 3840
rect 2650 3836 2654 3840
rect 2672 3836 2676 3840
rect 2680 3836 2684 3840
rect 2745 3836 2749 3840
rect 2817 3836 2821 3840
rect 2825 3836 2829 3840
rect 2897 3836 2901 3840
rect 2905 3836 2909 3840
rect 2977 3836 2981 3840
rect 2985 3836 2989 3840
rect 3031 3836 3035 3840
rect 3105 3836 3109 3840
rect 3156 3836 3160 3840
rect 3164 3836 3168 3840
rect 3186 3836 3190 3840
rect 3265 3836 3269 3840
rect 3285 3836 3289 3840
rect 3305 3836 3309 3840
rect 3351 3836 3355 3840
rect 3371 3836 3375 3840
rect 3391 3836 3395 3840
rect 3451 3836 3455 3840
rect 3511 3836 3515 3840
rect 3533 3836 3537 3840
rect 3555 3836 3559 3840
rect 3616 3836 3620 3840
rect 3624 3836 3628 3840
rect 3646 3836 3650 3840
rect 3716 3836 3720 3840
rect 3724 3836 3728 3840
rect 3746 3836 3750 3840
rect 3815 3836 3819 3840
rect 3835 3836 3839 3840
rect 3849 3836 3853 3840
rect 3869 3836 3873 3840
rect 3881 3836 3885 3840
rect 3901 3836 3905 3840
rect 3947 3836 3951 3840
rect 3955 3836 3959 3840
rect 3975 3836 3979 3840
rect 3983 3836 3987 3840
rect 4005 3836 4009 3840
rect 4051 3836 4055 3840
rect 4073 3836 4077 3840
rect 4157 3836 4161 3840
rect 4165 3836 4169 3840
rect 4211 3836 4215 3840
rect 4231 3836 4235 3840
rect 4251 3836 4255 3840
rect 4311 3836 4315 3840
rect 4333 3836 4337 3840
rect 4341 3836 4345 3840
rect 4361 3836 4365 3840
rect 4369 3836 4373 3840
rect 4415 3836 4419 3840
rect 4435 3836 4439 3840
rect 4447 3836 4451 3840
rect 4467 3836 4471 3840
rect 4481 3836 4485 3840
rect 4501 3836 4505 3840
rect 4551 3836 4555 3840
rect 4573 3836 4577 3840
rect 4645 3836 4649 3840
rect 4691 3836 4695 3840
rect 57 3733 61 3756
rect 46 3721 61 3733
rect 65 3733 69 3756
rect 116 3752 120 3756
rect 102 3744 120 3752
rect 102 3733 106 3744
rect 65 3721 74 3733
rect 45 3644 49 3721
rect 65 3644 69 3721
rect 102 3676 106 3721
rect 124 3699 128 3756
rect 146 3753 150 3796
rect 146 3741 153 3753
rect 126 3687 135 3699
rect 102 3669 115 3676
rect 111 3664 115 3669
rect 131 3664 135 3687
rect 151 3664 155 3741
rect 225 3713 229 3796
rect 225 3701 234 3713
rect 225 3644 229 3701
rect 285 3699 289 3756
rect 305 3742 309 3756
rect 325 3742 329 3756
rect 305 3736 320 3742
rect 325 3736 341 3742
rect 314 3713 320 3736
rect 285 3687 294 3699
rect 292 3644 296 3687
rect 314 3664 318 3701
rect 334 3699 341 3736
rect 334 3674 341 3687
rect 322 3668 341 3674
rect 381 3682 385 3756
rect 403 3719 407 3796
rect 425 3733 429 3796
rect 425 3721 434 3733
rect 406 3707 419 3719
rect 381 3670 393 3682
rect 322 3664 326 3668
rect 395 3664 399 3670
rect 415 3664 419 3707
rect 425 3664 429 3721
rect 485 3719 489 3796
rect 486 3707 489 3719
rect 483 3691 489 3707
rect 505 3719 509 3796
rect 565 3719 569 3796
rect 505 3707 514 3719
rect 566 3707 569 3719
rect 505 3691 511 3707
rect 483 3684 497 3691
rect 493 3664 497 3684
rect 503 3684 511 3691
rect 563 3691 569 3707
rect 585 3719 589 3796
rect 585 3707 594 3719
rect 631 3713 635 3796
rect 696 3752 700 3756
rect 682 3744 700 3752
rect 682 3733 686 3744
rect 585 3691 591 3707
rect 626 3701 635 3713
rect 563 3684 577 3691
rect 503 3664 507 3684
rect 573 3664 577 3684
rect 583 3684 591 3691
rect 583 3664 587 3684
rect 631 3644 635 3701
rect 682 3676 686 3721
rect 704 3699 708 3756
rect 726 3753 730 3796
rect 726 3741 733 3753
rect 706 3687 715 3699
rect 682 3669 695 3676
rect 691 3664 695 3669
rect 711 3664 715 3687
rect 731 3664 735 3741
rect 791 3719 795 3796
rect 786 3707 795 3719
rect 789 3691 795 3707
rect 811 3719 815 3796
rect 885 3753 889 3796
rect 905 3784 909 3796
rect 925 3788 929 3796
rect 925 3784 940 3788
rect 905 3780 920 3784
rect 914 3773 920 3780
rect 885 3741 893 3753
rect 905 3741 912 3753
rect 811 3707 814 3719
rect 811 3691 817 3707
rect 789 3684 797 3691
rect 793 3664 797 3684
rect 803 3684 817 3691
rect 908 3684 912 3741
rect 916 3684 920 3761
rect 934 3753 940 3784
rect 1071 3788 1075 3796
rect 1060 3784 1075 3788
rect 1091 3784 1095 3796
rect 924 3741 934 3753
rect 971 3742 975 3756
rect 991 3742 995 3756
rect 924 3684 928 3741
rect 959 3736 975 3742
rect 980 3736 995 3742
rect 959 3699 966 3736
rect 980 3713 986 3736
rect 803 3664 807 3684
rect 959 3674 966 3687
rect 959 3668 978 3674
rect 974 3664 978 3668
rect 982 3664 986 3701
rect 1011 3699 1015 3756
rect 1060 3753 1066 3784
rect 1080 3780 1095 3784
rect 1080 3773 1086 3780
rect 1066 3741 1076 3753
rect 1006 3687 1015 3699
rect 1004 3644 1008 3687
rect 1072 3684 1076 3741
rect 1080 3684 1084 3761
rect 1111 3753 1115 3796
rect 1088 3741 1095 3753
rect 1107 3741 1115 3753
rect 1171 3742 1175 3756
rect 1191 3742 1195 3756
rect 1088 3684 1092 3741
rect 1159 3736 1175 3742
rect 1180 3736 1195 3742
rect 1159 3699 1166 3736
rect 1180 3713 1186 3736
rect 1159 3674 1166 3687
rect 1159 3668 1178 3674
rect 1174 3664 1178 3668
rect 1182 3664 1186 3701
rect 1211 3699 1215 3756
rect 1271 3713 1275 3796
rect 1345 3753 1349 3796
rect 1365 3784 1369 3796
rect 1385 3788 1389 3796
rect 1385 3784 1400 3788
rect 1365 3780 1380 3784
rect 1374 3773 1380 3780
rect 1345 3741 1353 3753
rect 1365 3741 1372 3753
rect 1266 3701 1275 3713
rect 1206 3687 1215 3699
rect 1204 3644 1208 3687
rect 1271 3644 1275 3701
rect 1368 3684 1372 3741
rect 1376 3684 1380 3761
rect 1394 3753 1400 3784
rect 1384 3741 1394 3753
rect 1384 3684 1388 3741
rect 1445 3713 1449 3796
rect 1510 3753 1514 3796
rect 1507 3741 1514 3753
rect 1445 3701 1454 3713
rect 1445 3644 1449 3701
rect 1505 3664 1509 3741
rect 1532 3699 1536 3756
rect 1540 3752 1544 3756
rect 1540 3744 1558 3752
rect 1554 3733 1558 3744
rect 1525 3687 1534 3699
rect 1525 3664 1529 3687
rect 1554 3676 1558 3721
rect 1545 3669 1558 3676
rect 1605 3713 1609 3796
rect 1651 3742 1655 3756
rect 1671 3742 1675 3756
rect 1639 3736 1655 3742
rect 1660 3736 1675 3742
rect 1605 3701 1614 3713
rect 1545 3664 1549 3669
rect 1605 3644 1609 3701
rect 1639 3699 1646 3736
rect 1660 3713 1666 3736
rect 1639 3674 1646 3687
rect 1639 3668 1658 3674
rect 1654 3664 1658 3668
rect 1662 3664 1666 3701
rect 1691 3699 1695 3756
rect 1751 3733 1755 3756
rect 1746 3721 1755 3733
rect 1759 3733 1763 3756
rect 1759 3721 1774 3733
rect 1686 3687 1695 3699
rect 1684 3644 1688 3687
rect 1751 3644 1755 3721
rect 1771 3644 1775 3721
rect 1845 3699 1849 3756
rect 1865 3742 1869 3756
rect 1885 3742 1889 3756
rect 1865 3736 1880 3742
rect 1885 3736 1901 3742
rect 1874 3713 1880 3736
rect 1845 3687 1854 3699
rect 1852 3644 1856 3687
rect 1874 3664 1878 3701
rect 1894 3699 1901 3736
rect 1945 3719 1949 3796
rect 1946 3707 1949 3719
rect 1943 3691 1949 3707
rect 1965 3719 1969 3796
rect 2011 3752 2015 3756
rect 2002 3747 2015 3752
rect 1965 3707 1974 3719
rect 2002 3713 2006 3747
rect 2021 3733 2025 3756
rect 2041 3751 2045 3756
rect 2111 3733 2115 3796
rect 2133 3750 2137 3756
rect 2135 3738 2137 3750
rect 2106 3721 2115 3733
rect 1965 3691 1971 3707
rect 1894 3674 1901 3687
rect 1943 3684 1957 3691
rect 1882 3668 1901 3674
rect 1882 3664 1886 3668
rect 1953 3664 1957 3684
rect 1963 3684 1971 3691
rect 1963 3664 1967 3684
rect 2002 3656 2006 3701
rect 2021 3657 2025 3721
rect 2045 3672 2055 3684
rect 2051 3664 2055 3672
rect 2002 3651 2015 3656
rect 2021 3651 2035 3657
rect 2011 3644 2015 3651
rect 2031 3644 2035 3651
rect 2111 3644 2115 3721
rect 2205 3696 2209 3756
rect 2225 3696 2229 3756
rect 2245 3696 2249 3756
rect 2265 3696 2269 3756
rect 2285 3696 2289 3756
rect 2305 3696 2309 3756
rect 2325 3699 2329 3756
rect 2345 3699 2349 3756
rect 2395 3713 2399 3756
rect 2415 3714 2419 3796
rect 2429 3737 2433 3796
rect 2449 3756 2453 3796
rect 2461 3790 2465 3796
rect 2455 3744 2458 3756
rect 2429 3729 2438 3737
rect 2205 3684 2218 3696
rect 2245 3684 2258 3696
rect 2285 3684 2298 3696
rect 2325 3687 2334 3699
rect 2346 3687 2349 3699
rect 2135 3670 2137 3682
rect 2133 3664 2137 3670
rect 2205 3664 2209 3684
rect 2225 3664 2229 3684
rect 2245 3664 2249 3684
rect 2265 3664 2269 3684
rect 2285 3664 2289 3684
rect 2305 3664 2309 3684
rect 2325 3664 2329 3687
rect 2345 3664 2349 3687
rect 2395 3664 2399 3701
rect 2415 3644 2419 3702
rect 2434 3700 2438 3729
rect 2454 3680 2458 3744
rect 2425 3676 2458 3680
rect 2425 3644 2429 3676
rect 2463 3668 2467 3778
rect 2481 3770 2485 3796
rect 2527 3792 2531 3796
rect 2495 3790 2531 3792
rect 2507 3788 2531 3790
rect 2449 3656 2451 3668
rect 2447 3644 2451 3656
rect 2457 3656 2459 3668
rect 2457 3644 2461 3656
rect 2479 3644 2483 3758
rect 2495 3652 2499 3778
rect 2535 3764 2539 3796
rect 2555 3776 2559 3816
rect 2563 3793 2567 3816
rect 2563 3786 2571 3793
rect 2533 3669 2539 3764
rect 2567 3757 2571 3786
rect 2563 3751 2571 3757
rect 2563 3705 2567 3751
rect 2585 3744 2589 3756
rect 2650 3753 2654 3796
rect 2587 3732 2589 3744
rect 2647 3741 2654 3753
rect 2533 3665 2557 3669
rect 2519 3660 2537 3661
rect 2507 3656 2537 3660
rect 2495 3648 2529 3652
rect 2525 3644 2529 3648
rect 2533 3644 2537 3656
rect 2553 3644 2557 3665
rect 2563 3644 2567 3693
rect 2585 3664 2589 3732
rect 2645 3664 2649 3741
rect 2672 3699 2676 3756
rect 2680 3752 2684 3756
rect 2680 3744 2698 3752
rect 2694 3733 2698 3744
rect 2665 3687 2674 3699
rect 2665 3664 2669 3687
rect 2694 3676 2698 3721
rect 2685 3669 2698 3676
rect 2745 3713 2749 3796
rect 2817 3733 2821 3756
rect 2806 3721 2821 3733
rect 2825 3733 2829 3756
rect 2897 3733 2901 3756
rect 2825 3721 2834 3733
rect 2886 3721 2901 3733
rect 2905 3733 2909 3756
rect 2977 3733 2981 3756
rect 2905 3721 2914 3733
rect 2966 3721 2981 3733
rect 2985 3733 2989 3756
rect 2985 3721 2994 3733
rect 2745 3701 2754 3713
rect 2685 3664 2689 3669
rect 2745 3644 2749 3701
rect 2805 3644 2809 3721
rect 2825 3644 2829 3721
rect 2885 3644 2889 3721
rect 2905 3644 2909 3721
rect 2965 3644 2969 3721
rect 2985 3644 2989 3721
rect 3031 3713 3035 3796
rect 3026 3701 3035 3713
rect 3031 3644 3035 3701
rect 3105 3713 3109 3796
rect 3156 3752 3160 3756
rect 3142 3744 3160 3752
rect 3142 3733 3146 3744
rect 3105 3701 3114 3713
rect 3105 3644 3109 3701
rect 3142 3676 3146 3721
rect 3164 3699 3168 3756
rect 3186 3753 3190 3796
rect 3186 3741 3193 3753
rect 3166 3687 3175 3699
rect 3142 3669 3155 3676
rect 3151 3664 3155 3669
rect 3171 3664 3175 3687
rect 3191 3664 3195 3741
rect 3265 3699 3269 3756
rect 3285 3742 3289 3756
rect 3305 3742 3309 3756
rect 3351 3742 3355 3756
rect 3371 3742 3375 3756
rect 3285 3736 3300 3742
rect 3305 3736 3321 3742
rect 3294 3713 3300 3736
rect 3265 3687 3274 3699
rect 3272 3644 3276 3687
rect 3294 3664 3298 3701
rect 3314 3699 3321 3736
rect 3339 3736 3355 3742
rect 3360 3736 3375 3742
rect 3339 3699 3346 3736
rect 3360 3713 3366 3736
rect 3314 3674 3321 3687
rect 3302 3668 3321 3674
rect 3339 3674 3346 3687
rect 3339 3668 3358 3674
rect 3302 3664 3306 3668
rect 3354 3664 3358 3668
rect 3362 3664 3366 3701
rect 3391 3699 3395 3756
rect 3451 3713 3455 3796
rect 3511 3733 3515 3796
rect 3506 3721 3515 3733
rect 3446 3701 3455 3713
rect 3386 3687 3395 3699
rect 3384 3644 3388 3687
rect 3451 3644 3455 3701
rect 3511 3664 3515 3721
rect 3533 3719 3537 3796
rect 3521 3707 3534 3719
rect 3521 3664 3525 3707
rect 3555 3682 3559 3756
rect 3616 3752 3620 3756
rect 3602 3744 3620 3752
rect 3602 3733 3606 3744
rect 3547 3670 3559 3682
rect 3602 3676 3606 3721
rect 3624 3699 3628 3756
rect 3646 3753 3650 3796
rect 3646 3741 3653 3753
rect 3716 3752 3720 3756
rect 3702 3744 3720 3752
rect 3626 3687 3635 3699
rect 3541 3664 3545 3670
rect 3602 3669 3615 3676
rect 3611 3664 3615 3669
rect 3631 3664 3635 3687
rect 3651 3664 3655 3741
rect 3702 3733 3706 3744
rect 3702 3676 3706 3721
rect 3724 3699 3728 3756
rect 3746 3753 3750 3796
rect 3746 3741 3753 3753
rect 3726 3687 3735 3699
rect 3702 3669 3715 3676
rect 3711 3664 3715 3669
rect 3731 3664 3735 3687
rect 3751 3664 3755 3741
rect 3815 3713 3819 3756
rect 3835 3714 3839 3796
rect 3849 3737 3853 3796
rect 3869 3756 3873 3796
rect 3881 3790 3885 3796
rect 3875 3744 3878 3756
rect 3849 3729 3858 3737
rect 3815 3664 3819 3701
rect 3835 3644 3839 3702
rect 3854 3700 3858 3729
rect 3874 3680 3878 3744
rect 3845 3676 3878 3680
rect 3845 3644 3849 3676
rect 3883 3668 3887 3778
rect 3901 3770 3905 3796
rect 3947 3792 3951 3796
rect 3915 3790 3951 3792
rect 3927 3788 3951 3790
rect 3869 3656 3871 3668
rect 3867 3644 3871 3656
rect 3877 3656 3879 3668
rect 3877 3644 3881 3656
rect 3899 3644 3903 3758
rect 3915 3652 3919 3778
rect 3955 3764 3959 3796
rect 3975 3776 3979 3816
rect 3983 3793 3987 3816
rect 3983 3786 3991 3793
rect 3953 3669 3959 3764
rect 3987 3757 3991 3786
rect 3983 3751 3991 3757
rect 3983 3705 3987 3751
rect 4005 3744 4009 3756
rect 4007 3732 4009 3744
rect 4051 3733 4055 3796
rect 4333 3793 4337 3816
rect 4329 3786 4337 3793
rect 4329 3757 4333 3786
rect 4341 3776 4345 3816
rect 4361 3764 4365 3796
rect 4369 3792 4373 3796
rect 4369 3790 4405 3792
rect 4369 3788 4393 3790
rect 4073 3750 4077 3756
rect 4075 3738 4077 3750
rect 4157 3733 4161 3756
rect 3953 3665 3977 3669
rect 3939 3660 3957 3661
rect 3927 3656 3957 3660
rect 3915 3648 3949 3652
rect 3945 3644 3949 3648
rect 3953 3644 3957 3656
rect 3973 3644 3977 3665
rect 3983 3644 3987 3693
rect 4005 3664 4009 3732
rect 4046 3721 4055 3733
rect 4146 3721 4161 3733
rect 4165 3733 4169 3756
rect 4211 3742 4215 3756
rect 4231 3742 4235 3756
rect 4199 3736 4215 3742
rect 4220 3736 4235 3742
rect 4165 3721 4174 3733
rect 4051 3644 4055 3721
rect 4075 3670 4077 3682
rect 4073 3664 4077 3670
rect 4145 3644 4149 3721
rect 4165 3644 4169 3721
rect 4199 3699 4206 3736
rect 4220 3713 4226 3736
rect 4199 3674 4206 3687
rect 4199 3668 4218 3674
rect 4214 3664 4218 3668
rect 4222 3664 4226 3701
rect 4251 3699 4255 3756
rect 4246 3687 4255 3699
rect 4311 3744 4315 3756
rect 4329 3751 4337 3757
rect 4311 3732 4313 3744
rect 4244 3644 4248 3687
rect 4311 3664 4315 3732
rect 4333 3705 4337 3751
rect 4333 3644 4337 3693
rect 4361 3669 4367 3764
rect 4343 3665 4367 3669
rect 4343 3644 4347 3665
rect 4363 3660 4381 3661
rect 4363 3656 4393 3660
rect 4363 3644 4367 3656
rect 4401 3652 4405 3778
rect 4415 3770 4419 3796
rect 4435 3790 4439 3796
rect 4371 3648 4405 3652
rect 4371 3644 4375 3648
rect 4417 3644 4421 3758
rect 4433 3668 4437 3778
rect 4447 3756 4451 3796
rect 4442 3744 4445 3756
rect 4442 3680 4446 3744
rect 4467 3737 4471 3796
rect 4462 3729 4471 3737
rect 4462 3700 4466 3729
rect 4481 3714 4485 3796
rect 4501 3713 4505 3756
rect 4551 3733 4555 3796
rect 4573 3750 4577 3756
rect 4575 3738 4577 3750
rect 4546 3721 4555 3733
rect 4442 3676 4475 3680
rect 4441 3656 4443 3668
rect 4439 3644 4443 3656
rect 4449 3656 4451 3668
rect 4449 3644 4453 3656
rect 4471 3644 4475 3676
rect 4481 3644 4485 3702
rect 4501 3664 4505 3701
rect 4551 3644 4555 3721
rect 4645 3713 4649 3796
rect 4691 3713 4695 3796
rect 4645 3701 4654 3713
rect 4686 3701 4695 3713
rect 4575 3670 4577 3682
rect 4573 3664 4577 3670
rect 4645 3644 4649 3701
rect 4691 3644 4695 3701
rect 45 3620 49 3624
rect 65 3620 69 3624
rect 111 3620 115 3624
rect 131 3620 135 3624
rect 151 3620 155 3624
rect 225 3620 229 3624
rect 292 3620 296 3624
rect 314 3620 318 3624
rect 322 3620 326 3624
rect 395 3620 399 3624
rect 415 3620 419 3624
rect 425 3620 429 3624
rect 493 3620 497 3624
rect 503 3620 507 3624
rect 573 3620 577 3624
rect 583 3620 587 3624
rect 631 3620 635 3624
rect 691 3620 695 3624
rect 711 3620 715 3624
rect 731 3620 735 3624
rect 793 3620 797 3624
rect 803 3620 807 3624
rect 908 3620 912 3624
rect 916 3620 920 3624
rect 924 3620 928 3624
rect 974 3620 978 3624
rect 982 3620 986 3624
rect 1004 3620 1008 3624
rect 1072 3620 1076 3624
rect 1080 3620 1084 3624
rect 1088 3620 1092 3624
rect 1174 3620 1178 3624
rect 1182 3620 1186 3624
rect 1204 3620 1208 3624
rect 1271 3620 1275 3624
rect 1368 3620 1372 3624
rect 1376 3620 1380 3624
rect 1384 3620 1388 3624
rect 1445 3620 1449 3624
rect 1505 3620 1509 3624
rect 1525 3620 1529 3624
rect 1545 3620 1549 3624
rect 1605 3620 1609 3624
rect 1654 3620 1658 3624
rect 1662 3620 1666 3624
rect 1684 3620 1688 3624
rect 1751 3620 1755 3624
rect 1771 3620 1775 3624
rect 1852 3620 1856 3624
rect 1874 3620 1878 3624
rect 1882 3620 1886 3624
rect 1953 3620 1957 3624
rect 1963 3620 1967 3624
rect 2011 3620 2015 3624
rect 2031 3620 2035 3624
rect 2051 3620 2055 3624
rect 2111 3620 2115 3624
rect 2133 3620 2137 3624
rect 2205 3620 2209 3624
rect 2225 3620 2229 3624
rect 2245 3620 2249 3624
rect 2265 3620 2269 3624
rect 2285 3620 2289 3624
rect 2305 3620 2309 3624
rect 2325 3620 2329 3624
rect 2345 3620 2349 3624
rect 2395 3620 2399 3624
rect 2415 3620 2419 3624
rect 2425 3620 2429 3624
rect 2447 3620 2451 3624
rect 2457 3620 2461 3624
rect 2479 3620 2483 3624
rect 2525 3620 2529 3624
rect 2533 3620 2537 3624
rect 2553 3620 2557 3624
rect 2563 3620 2567 3624
rect 2585 3620 2589 3624
rect 2645 3620 2649 3624
rect 2665 3620 2669 3624
rect 2685 3620 2689 3624
rect 2745 3620 2749 3624
rect 2805 3620 2809 3624
rect 2825 3620 2829 3624
rect 2885 3620 2889 3624
rect 2905 3620 2909 3624
rect 2965 3620 2969 3624
rect 2985 3620 2989 3624
rect 3031 3620 3035 3624
rect 3105 3620 3109 3624
rect 3151 3620 3155 3624
rect 3171 3620 3175 3624
rect 3191 3620 3195 3624
rect 3272 3620 3276 3624
rect 3294 3620 3298 3624
rect 3302 3620 3306 3624
rect 3354 3620 3358 3624
rect 3362 3620 3366 3624
rect 3384 3620 3388 3624
rect 3451 3620 3455 3624
rect 3511 3620 3515 3624
rect 3521 3620 3525 3624
rect 3541 3620 3545 3624
rect 3611 3620 3615 3624
rect 3631 3620 3635 3624
rect 3651 3620 3655 3624
rect 3711 3620 3715 3624
rect 3731 3620 3735 3624
rect 3751 3620 3755 3624
rect 3815 3620 3819 3624
rect 3835 3620 3839 3624
rect 3845 3620 3849 3624
rect 3867 3620 3871 3624
rect 3877 3620 3881 3624
rect 3899 3620 3903 3624
rect 3945 3620 3949 3624
rect 3953 3620 3957 3624
rect 3973 3620 3977 3624
rect 3983 3620 3987 3624
rect 4005 3620 4009 3624
rect 4051 3620 4055 3624
rect 4073 3620 4077 3624
rect 4145 3620 4149 3624
rect 4165 3620 4169 3624
rect 4214 3620 4218 3624
rect 4222 3620 4226 3624
rect 4244 3620 4248 3624
rect 4311 3620 4315 3624
rect 4333 3620 4337 3624
rect 4343 3620 4347 3624
rect 4363 3620 4367 3624
rect 4371 3620 4375 3624
rect 4417 3620 4421 3624
rect 4439 3620 4443 3624
rect 4449 3620 4453 3624
rect 4471 3620 4475 3624
rect 4481 3620 4485 3624
rect 4501 3620 4505 3624
rect 4551 3620 4555 3624
rect 4573 3620 4577 3624
rect 4645 3620 4649 3624
rect 4691 3620 4695 3624
rect 53 3596 57 3600
rect 63 3596 67 3600
rect 115 3596 119 3600
rect 135 3596 139 3600
rect 145 3596 149 3600
rect 167 3596 171 3600
rect 177 3596 181 3600
rect 199 3596 203 3600
rect 245 3596 249 3600
rect 253 3596 257 3600
rect 273 3596 277 3600
rect 283 3596 287 3600
rect 305 3596 309 3600
rect 365 3596 369 3600
rect 433 3596 437 3600
rect 443 3596 447 3600
rect 505 3596 509 3600
rect 525 3596 529 3600
rect 545 3596 549 3600
rect 605 3596 609 3600
rect 625 3596 629 3600
rect 645 3596 649 3600
rect 693 3596 697 3600
rect 703 3596 707 3600
rect 771 3596 775 3600
rect 791 3596 795 3600
rect 811 3596 815 3600
rect 831 3596 835 3600
rect 891 3596 895 3600
rect 988 3596 992 3600
rect 996 3596 1000 3600
rect 1004 3596 1008 3600
rect 1054 3596 1058 3600
rect 1062 3596 1066 3600
rect 1084 3596 1088 3600
rect 1151 3596 1155 3600
rect 1171 3596 1175 3600
rect 1233 3596 1237 3600
rect 1243 3596 1247 3600
rect 1313 3596 1317 3600
rect 1323 3596 1327 3600
rect 1391 3596 1395 3600
rect 1411 3596 1415 3600
rect 1431 3596 1435 3600
rect 1495 3596 1499 3600
rect 1515 3596 1519 3600
rect 1525 3596 1529 3600
rect 1547 3596 1551 3600
rect 1557 3596 1561 3600
rect 1579 3596 1583 3600
rect 1625 3596 1629 3600
rect 1633 3596 1637 3600
rect 1653 3596 1657 3600
rect 1663 3596 1667 3600
rect 1685 3596 1689 3600
rect 1753 3596 1757 3600
rect 1763 3596 1767 3600
rect 1811 3596 1815 3600
rect 1831 3596 1835 3600
rect 1851 3596 1855 3600
rect 1911 3596 1915 3600
rect 1993 3596 1997 3600
rect 2003 3596 2007 3600
rect 2075 3596 2079 3600
rect 2095 3596 2099 3600
rect 2105 3596 2109 3600
rect 2153 3596 2157 3600
rect 2163 3596 2167 3600
rect 2232 3596 2236 3600
rect 2240 3596 2244 3600
rect 2248 3596 2252 3600
rect 2331 3596 2335 3600
rect 2391 3596 2395 3600
rect 2451 3596 2455 3600
rect 2473 3596 2477 3600
rect 2483 3596 2487 3600
rect 2503 3596 2507 3600
rect 2511 3596 2515 3600
rect 2557 3596 2561 3600
rect 2579 3596 2583 3600
rect 2589 3596 2593 3600
rect 2611 3596 2615 3600
rect 2621 3596 2625 3600
rect 2641 3596 2645 3600
rect 2691 3596 2695 3600
rect 2711 3596 2715 3600
rect 2731 3596 2735 3600
rect 2791 3596 2795 3600
rect 2813 3596 2817 3600
rect 2873 3596 2877 3600
rect 2883 3596 2887 3600
rect 2951 3596 2955 3600
rect 2973 3596 2977 3600
rect 2983 3596 2987 3600
rect 3003 3596 3007 3600
rect 3011 3596 3015 3600
rect 3057 3596 3061 3600
rect 3079 3596 3083 3600
rect 3089 3596 3093 3600
rect 3111 3596 3115 3600
rect 3121 3596 3125 3600
rect 3141 3596 3145 3600
rect 3205 3596 3209 3600
rect 3225 3596 3229 3600
rect 3245 3596 3249 3600
rect 3305 3596 3309 3600
rect 3351 3596 3355 3600
rect 3371 3596 3375 3600
rect 3431 3596 3435 3600
rect 3505 3596 3509 3600
rect 3525 3596 3529 3600
rect 3574 3596 3578 3600
rect 3582 3596 3586 3600
rect 3604 3596 3608 3600
rect 3671 3596 3675 3600
rect 3691 3596 3695 3600
rect 3711 3596 3715 3600
rect 3806 3596 3810 3600
rect 3814 3596 3818 3600
rect 3834 3596 3838 3600
rect 3842 3596 3846 3600
rect 3913 3596 3917 3600
rect 3923 3596 3927 3600
rect 3971 3596 3975 3600
rect 3993 3596 3997 3600
rect 4003 3596 4007 3600
rect 4023 3596 4027 3600
rect 4031 3596 4035 3600
rect 4077 3596 4081 3600
rect 4099 3596 4103 3600
rect 4109 3596 4113 3600
rect 4131 3596 4135 3600
rect 4141 3596 4145 3600
rect 4161 3596 4165 3600
rect 4211 3596 4215 3600
rect 4233 3596 4237 3600
rect 4243 3596 4247 3600
rect 4263 3596 4267 3600
rect 4271 3596 4275 3600
rect 4317 3596 4321 3600
rect 4339 3596 4343 3600
rect 4349 3596 4353 3600
rect 4371 3596 4375 3600
rect 4381 3596 4385 3600
rect 4401 3596 4405 3600
rect 4465 3596 4469 3600
rect 4485 3596 4489 3600
rect 4505 3596 4509 3600
rect 4525 3596 4529 3600
rect 4545 3596 4549 3600
rect 4565 3596 4569 3600
rect 4585 3596 4589 3600
rect 4605 3596 4609 3600
rect 4651 3596 4655 3600
rect 4671 3596 4675 3600
rect 4691 3596 4695 3600
rect 53 3536 57 3556
rect 43 3529 57 3536
rect 63 3536 67 3556
rect 63 3529 71 3536
rect 43 3513 49 3529
rect 46 3501 49 3513
rect 45 3424 49 3501
rect 65 3513 71 3529
rect 115 3519 119 3556
rect 65 3501 74 3513
rect 135 3518 139 3576
rect 145 3544 149 3576
rect 167 3564 171 3576
rect 169 3552 171 3564
rect 177 3564 181 3576
rect 177 3552 179 3564
rect 145 3540 178 3544
rect 65 3424 69 3501
rect 115 3464 119 3507
rect 135 3424 139 3506
rect 154 3491 158 3520
rect 149 3483 158 3491
rect 149 3424 153 3483
rect 174 3476 178 3540
rect 175 3464 178 3476
rect 169 3424 173 3464
rect 183 3442 187 3552
rect 199 3462 203 3576
rect 245 3572 249 3576
rect 215 3568 249 3572
rect 181 3424 185 3430
rect 201 3424 205 3450
rect 215 3442 219 3568
rect 253 3564 257 3576
rect 227 3560 257 3564
rect 239 3559 257 3560
rect 273 3555 277 3576
rect 253 3551 277 3555
rect 253 3456 259 3551
rect 283 3527 287 3576
rect 283 3469 287 3515
rect 305 3488 309 3556
rect 307 3476 309 3488
rect 283 3463 291 3469
rect 305 3464 309 3476
rect 365 3519 369 3576
rect 433 3536 437 3556
rect 423 3529 437 3536
rect 443 3536 447 3556
rect 443 3529 451 3536
rect 365 3507 374 3519
rect 423 3513 429 3529
rect 227 3430 251 3432
rect 215 3428 251 3430
rect 247 3424 251 3428
rect 255 3424 259 3456
rect 275 3404 279 3444
rect 287 3434 291 3463
rect 283 3427 291 3434
rect 283 3404 287 3427
rect 365 3424 369 3507
rect 426 3501 429 3513
rect 425 3424 429 3501
rect 445 3513 451 3529
rect 445 3501 454 3513
rect 445 3424 449 3501
rect 505 3479 509 3556
rect 525 3533 529 3556
rect 545 3551 549 3556
rect 545 3544 558 3551
rect 525 3521 534 3533
rect 507 3467 514 3479
rect 510 3424 514 3467
rect 532 3464 536 3521
rect 554 3499 558 3544
rect 554 3476 558 3487
rect 605 3479 609 3556
rect 625 3533 629 3556
rect 645 3551 649 3556
rect 645 3544 658 3551
rect 625 3521 634 3533
rect 540 3468 558 3476
rect 540 3464 544 3468
rect 607 3467 614 3479
rect 610 3424 614 3467
rect 632 3464 636 3521
rect 654 3499 658 3544
rect 693 3536 697 3556
rect 689 3529 697 3536
rect 703 3536 707 3556
rect 771 3549 775 3556
rect 760 3545 775 3549
rect 703 3529 717 3536
rect 689 3513 695 3529
rect 686 3501 695 3513
rect 654 3476 658 3487
rect 640 3468 658 3476
rect 640 3464 644 3468
rect 691 3424 695 3501
rect 711 3513 717 3529
rect 711 3501 714 3513
rect 711 3424 715 3501
rect 760 3499 766 3545
rect 791 3533 795 3556
rect 811 3533 815 3556
rect 786 3521 795 3533
rect 761 3472 766 3487
rect 789 3472 795 3521
rect 761 3468 775 3472
rect 771 3464 775 3468
rect 781 3468 795 3472
rect 781 3464 785 3468
rect 811 3464 815 3521
rect 831 3499 835 3556
rect 891 3519 895 3576
rect 1054 3552 1058 3556
rect 1039 3546 1058 3552
rect 886 3507 895 3519
rect 831 3487 833 3499
rect 831 3472 835 3487
rect 821 3468 835 3472
rect 821 3464 825 3468
rect 891 3424 895 3507
rect 988 3479 992 3536
rect 965 3467 973 3479
rect 985 3467 992 3479
rect 965 3424 969 3467
rect 996 3459 1000 3536
rect 1004 3479 1008 3536
rect 1039 3533 1046 3546
rect 1039 3484 1046 3521
rect 1062 3519 1066 3556
rect 1084 3533 1088 3576
rect 1086 3521 1095 3533
rect 1060 3484 1066 3507
rect 1004 3467 1014 3479
rect 1039 3478 1055 3484
rect 1060 3478 1075 3484
rect 994 3440 1000 3447
rect 985 3436 1000 3440
rect 1014 3436 1020 3467
rect 1051 3464 1055 3478
rect 1071 3464 1075 3478
rect 1091 3464 1095 3521
rect 1151 3499 1155 3576
rect 1171 3499 1175 3576
rect 1233 3536 1237 3556
rect 1229 3529 1237 3536
rect 1243 3536 1247 3556
rect 1313 3536 1317 3556
rect 1243 3529 1257 3536
rect 1229 3513 1235 3529
rect 1226 3501 1235 3513
rect 1146 3487 1155 3499
rect 1151 3464 1155 3487
rect 1159 3487 1174 3499
rect 1159 3464 1163 3487
rect 985 3424 989 3436
rect 1005 3432 1020 3436
rect 1005 3424 1009 3432
rect 1231 3424 1235 3501
rect 1251 3513 1257 3529
rect 1309 3529 1317 3536
rect 1323 3536 1327 3556
rect 1391 3551 1395 3556
rect 1382 3544 1395 3551
rect 1323 3529 1337 3536
rect 1309 3513 1315 3529
rect 1251 3501 1254 3513
rect 1306 3501 1315 3513
rect 1251 3424 1255 3501
rect 1311 3424 1315 3501
rect 1331 3513 1337 3529
rect 1331 3501 1334 3513
rect 1331 3424 1335 3501
rect 1382 3499 1386 3544
rect 1411 3533 1415 3556
rect 1406 3521 1415 3533
rect 1382 3476 1386 3487
rect 1382 3468 1400 3476
rect 1396 3464 1400 3468
rect 1404 3464 1408 3521
rect 1431 3479 1435 3556
rect 1495 3519 1499 3556
rect 1515 3518 1519 3576
rect 1525 3544 1529 3576
rect 1547 3564 1551 3576
rect 1549 3552 1551 3564
rect 1557 3564 1561 3576
rect 1557 3552 1559 3564
rect 1525 3540 1558 3544
rect 1426 3467 1433 3479
rect 1426 3424 1430 3467
rect 1495 3464 1499 3507
rect 1515 3424 1519 3506
rect 1534 3491 1538 3520
rect 1529 3483 1538 3491
rect 1529 3424 1533 3483
rect 1554 3476 1558 3540
rect 1555 3464 1558 3476
rect 1549 3424 1553 3464
rect 1563 3442 1567 3552
rect 1579 3462 1583 3576
rect 1625 3572 1629 3576
rect 1595 3568 1629 3572
rect 1561 3424 1565 3430
rect 1581 3424 1585 3450
rect 1595 3442 1599 3568
rect 1633 3564 1637 3576
rect 1607 3560 1637 3564
rect 1619 3559 1637 3560
rect 1653 3555 1657 3576
rect 1633 3551 1657 3555
rect 1633 3456 1639 3551
rect 1663 3527 1667 3576
rect 1663 3469 1667 3515
rect 1685 3488 1689 3556
rect 1753 3536 1757 3556
rect 1743 3529 1757 3536
rect 1763 3536 1767 3556
rect 1811 3551 1815 3556
rect 1802 3544 1815 3551
rect 1763 3529 1771 3536
rect 1743 3513 1749 3529
rect 1746 3501 1749 3513
rect 1687 3476 1689 3488
rect 1663 3463 1671 3469
rect 1685 3464 1689 3476
rect 1607 3430 1631 3432
rect 1595 3428 1631 3430
rect 1627 3424 1631 3428
rect 1635 3424 1639 3456
rect 1655 3404 1659 3444
rect 1667 3434 1671 3463
rect 1663 3427 1671 3434
rect 1663 3404 1667 3427
rect 1745 3424 1749 3501
rect 1765 3513 1771 3529
rect 1765 3501 1774 3513
rect 1765 3424 1769 3501
rect 1802 3499 1806 3544
rect 1831 3533 1835 3556
rect 1826 3521 1835 3533
rect 1802 3476 1806 3487
rect 1802 3468 1820 3476
rect 1816 3464 1820 3468
rect 1824 3464 1828 3521
rect 1851 3479 1855 3556
rect 1911 3533 1915 3556
rect 1993 3536 1997 3556
rect 1906 3521 1915 3533
rect 1846 3467 1853 3479
rect 1846 3424 1850 3467
rect 1911 3464 1915 3521
rect 1983 3529 1997 3536
rect 2003 3536 2007 3556
rect 2075 3550 2079 3556
rect 2061 3538 2073 3550
rect 2003 3529 2011 3536
rect 1983 3513 1989 3529
rect 1986 3501 1989 3513
rect 1985 3424 1989 3501
rect 2005 3513 2011 3529
rect 2005 3501 2014 3513
rect 2005 3424 2009 3501
rect 2061 3464 2065 3538
rect 2095 3513 2099 3556
rect 2086 3501 2099 3513
rect 2083 3424 2087 3501
rect 2105 3499 2109 3556
rect 2153 3536 2157 3556
rect 2149 3529 2157 3536
rect 2163 3536 2167 3556
rect 2163 3529 2177 3536
rect 2149 3513 2155 3529
rect 2146 3501 2155 3513
rect 2105 3487 2114 3499
rect 2105 3424 2109 3487
rect 2151 3424 2155 3501
rect 2171 3513 2177 3529
rect 2171 3501 2174 3513
rect 2171 3424 2175 3501
rect 2232 3479 2236 3536
rect 2226 3467 2236 3479
rect 2220 3436 2226 3467
rect 2240 3459 2244 3536
rect 2248 3479 2252 3536
rect 2331 3519 2335 3576
rect 2391 3519 2395 3576
rect 2326 3507 2335 3519
rect 2386 3507 2395 3519
rect 2248 3467 2255 3479
rect 2267 3467 2275 3479
rect 2240 3440 2246 3447
rect 2240 3436 2255 3440
rect 2220 3432 2235 3436
rect 2231 3424 2235 3432
rect 2251 3424 2255 3436
rect 2271 3424 2275 3467
rect 2331 3424 2335 3507
rect 2391 3424 2395 3507
rect 2451 3488 2455 3556
rect 2473 3527 2477 3576
rect 2483 3555 2487 3576
rect 2503 3564 2507 3576
rect 2511 3572 2515 3576
rect 2511 3568 2545 3572
rect 2503 3560 2533 3564
rect 2503 3559 2521 3560
rect 2483 3551 2507 3555
rect 2451 3476 2453 3488
rect 2451 3464 2455 3476
rect 2473 3469 2477 3515
rect 2469 3463 2477 3469
rect 2469 3434 2473 3463
rect 2501 3456 2507 3551
rect 2469 3427 2477 3434
rect 2473 3404 2477 3427
rect 2481 3404 2485 3444
rect 2501 3424 2505 3456
rect 2541 3442 2545 3568
rect 2557 3462 2561 3576
rect 2579 3564 2583 3576
rect 2581 3552 2583 3564
rect 2589 3564 2593 3576
rect 2589 3552 2591 3564
rect 2509 3430 2533 3432
rect 2509 3428 2545 3430
rect 2509 3424 2513 3428
rect 2555 3424 2559 3450
rect 2573 3442 2577 3552
rect 2611 3544 2615 3576
rect 2582 3540 2615 3544
rect 2582 3476 2586 3540
rect 2602 3491 2606 3520
rect 2621 3518 2625 3576
rect 2641 3519 2645 3556
rect 2691 3551 2695 3556
rect 2682 3544 2695 3551
rect 2602 3483 2611 3491
rect 2582 3464 2585 3476
rect 2575 3424 2579 3430
rect 2587 3424 2591 3464
rect 2607 3424 2611 3483
rect 2621 3424 2625 3506
rect 2641 3464 2645 3507
rect 2682 3499 2686 3544
rect 2711 3533 2715 3556
rect 2706 3521 2715 3533
rect 2682 3476 2686 3487
rect 2682 3468 2700 3476
rect 2696 3464 2700 3468
rect 2704 3464 2708 3521
rect 2731 3479 2735 3556
rect 2791 3499 2795 3576
rect 2813 3550 2817 3556
rect 2815 3538 2817 3550
rect 2873 3536 2877 3556
rect 2869 3529 2877 3536
rect 2883 3536 2887 3556
rect 2883 3529 2897 3536
rect 2869 3513 2875 3529
rect 2866 3501 2875 3513
rect 2786 3487 2795 3499
rect 2726 3467 2733 3479
rect 2726 3424 2730 3467
rect 2791 3424 2795 3487
rect 2815 3470 2817 3482
rect 2813 3464 2817 3470
rect 2871 3424 2875 3501
rect 2891 3513 2897 3529
rect 2891 3501 2894 3513
rect 2891 3424 2895 3501
rect 2951 3488 2955 3556
rect 2973 3527 2977 3576
rect 2983 3555 2987 3576
rect 3003 3564 3007 3576
rect 3011 3572 3015 3576
rect 3011 3568 3045 3572
rect 3003 3560 3033 3564
rect 3003 3559 3021 3560
rect 2983 3551 3007 3555
rect 2951 3476 2953 3488
rect 2951 3464 2955 3476
rect 2973 3469 2977 3515
rect 2969 3463 2977 3469
rect 2969 3434 2973 3463
rect 3001 3456 3007 3551
rect 2969 3427 2977 3434
rect 2973 3404 2977 3427
rect 2981 3404 2985 3444
rect 3001 3424 3005 3456
rect 3041 3442 3045 3568
rect 3057 3462 3061 3576
rect 3079 3564 3083 3576
rect 3081 3552 3083 3564
rect 3089 3564 3093 3576
rect 3089 3552 3091 3564
rect 3009 3430 3033 3432
rect 3009 3428 3045 3430
rect 3009 3424 3013 3428
rect 3055 3424 3059 3450
rect 3073 3442 3077 3552
rect 3111 3544 3115 3576
rect 3082 3540 3115 3544
rect 3082 3476 3086 3540
rect 3102 3491 3106 3520
rect 3121 3518 3125 3576
rect 3141 3519 3145 3556
rect 3102 3483 3111 3491
rect 3082 3464 3085 3476
rect 3075 3424 3079 3430
rect 3087 3424 3091 3464
rect 3107 3424 3111 3483
rect 3121 3424 3125 3506
rect 3141 3464 3145 3507
rect 3205 3479 3209 3556
rect 3225 3533 3229 3556
rect 3245 3551 3249 3556
rect 3245 3544 3258 3551
rect 3225 3521 3234 3533
rect 3207 3467 3214 3479
rect 3210 3424 3214 3467
rect 3232 3464 3236 3521
rect 3254 3499 3258 3544
rect 3305 3519 3309 3576
rect 3305 3507 3314 3519
rect 3254 3476 3258 3487
rect 3240 3468 3258 3476
rect 3240 3464 3244 3468
rect 3305 3424 3309 3507
rect 3351 3499 3355 3576
rect 3371 3499 3375 3576
rect 3431 3519 3435 3576
rect 3426 3507 3435 3519
rect 3346 3487 3355 3499
rect 3351 3464 3355 3487
rect 3359 3487 3374 3499
rect 3359 3464 3363 3487
rect 3431 3424 3435 3507
rect 3505 3499 3509 3576
rect 3525 3499 3529 3576
rect 3574 3552 3578 3556
rect 3559 3546 3578 3552
rect 3559 3533 3566 3546
rect 3506 3487 3521 3499
rect 3517 3464 3521 3487
rect 3525 3487 3534 3499
rect 3525 3464 3529 3487
rect 3559 3484 3566 3521
rect 3582 3519 3586 3556
rect 3604 3533 3608 3576
rect 3671 3569 3675 3576
rect 3691 3569 3695 3576
rect 3662 3564 3675 3569
rect 3606 3521 3615 3533
rect 3580 3484 3586 3507
rect 3559 3478 3575 3484
rect 3580 3478 3595 3484
rect 3571 3464 3575 3478
rect 3591 3464 3595 3478
rect 3611 3464 3615 3521
rect 3662 3519 3666 3564
rect 3662 3473 3666 3507
rect 3681 3563 3695 3569
rect 3681 3499 3685 3563
rect 3711 3548 3715 3556
rect 3806 3551 3810 3556
rect 3705 3536 3715 3548
rect 3780 3547 3810 3551
rect 3780 3499 3786 3547
rect 3814 3542 3818 3556
rect 3805 3535 3818 3542
rect 3805 3533 3809 3535
rect 3834 3533 3838 3556
rect 3842 3548 3846 3556
rect 3842 3541 3859 3548
rect 3807 3521 3809 3533
rect 3786 3487 3789 3499
rect 3662 3468 3675 3473
rect 3671 3464 3675 3468
rect 3681 3464 3685 3487
rect 3701 3464 3705 3469
rect 3785 3464 3789 3487
rect 3805 3464 3809 3521
rect 3834 3492 3838 3521
rect 3853 3499 3859 3541
rect 3913 3536 3917 3556
rect 3903 3529 3917 3536
rect 3923 3536 3927 3556
rect 3923 3529 3931 3536
rect 3903 3513 3909 3529
rect 3906 3501 3909 3513
rect 3825 3486 3838 3492
rect 3845 3487 3853 3492
rect 3845 3486 3865 3487
rect 3825 3464 3829 3486
rect 3845 3464 3849 3486
rect 3905 3424 3909 3501
rect 3925 3513 3931 3529
rect 3925 3501 3934 3513
rect 3925 3424 3929 3501
rect 3971 3488 3975 3556
rect 3993 3527 3997 3576
rect 4003 3555 4007 3576
rect 4023 3564 4027 3576
rect 4031 3572 4035 3576
rect 4031 3568 4065 3572
rect 4023 3560 4053 3564
rect 4023 3559 4041 3560
rect 4003 3551 4027 3555
rect 3971 3476 3973 3488
rect 3971 3464 3975 3476
rect 3993 3469 3997 3515
rect 3989 3463 3997 3469
rect 3989 3434 3993 3463
rect 4021 3456 4027 3551
rect 3989 3427 3997 3434
rect 3993 3404 3997 3427
rect 4001 3404 4005 3444
rect 4021 3424 4025 3456
rect 4061 3442 4065 3568
rect 4077 3462 4081 3576
rect 4099 3564 4103 3576
rect 4101 3552 4103 3564
rect 4109 3564 4113 3576
rect 4109 3552 4111 3564
rect 4029 3430 4053 3432
rect 4029 3428 4065 3430
rect 4029 3424 4033 3428
rect 4075 3424 4079 3450
rect 4093 3442 4097 3552
rect 4131 3544 4135 3576
rect 4102 3540 4135 3544
rect 4102 3476 4106 3540
rect 4122 3491 4126 3520
rect 4141 3518 4145 3576
rect 4161 3519 4165 3556
rect 4122 3483 4131 3491
rect 4102 3464 4105 3476
rect 4095 3424 4099 3430
rect 4107 3424 4111 3464
rect 4127 3424 4131 3483
rect 4141 3424 4145 3506
rect 4161 3464 4165 3507
rect 4211 3488 4215 3556
rect 4233 3527 4237 3576
rect 4243 3555 4247 3576
rect 4263 3564 4267 3576
rect 4271 3572 4275 3576
rect 4271 3568 4305 3572
rect 4263 3560 4293 3564
rect 4263 3559 4281 3560
rect 4243 3551 4267 3555
rect 4211 3476 4213 3488
rect 4211 3464 4215 3476
rect 4233 3469 4237 3515
rect 4229 3463 4237 3469
rect 4229 3434 4233 3463
rect 4261 3456 4267 3551
rect 4229 3427 4237 3434
rect 4233 3404 4237 3427
rect 4241 3404 4245 3444
rect 4261 3424 4265 3456
rect 4301 3442 4305 3568
rect 4317 3462 4321 3576
rect 4339 3564 4343 3576
rect 4341 3552 4343 3564
rect 4349 3564 4353 3576
rect 4349 3552 4351 3564
rect 4269 3430 4293 3432
rect 4269 3428 4305 3430
rect 4269 3424 4273 3428
rect 4315 3424 4319 3450
rect 4333 3442 4337 3552
rect 4371 3544 4375 3576
rect 4342 3540 4375 3544
rect 4342 3476 4346 3540
rect 4362 3491 4366 3520
rect 4381 3518 4385 3576
rect 4401 3519 4405 3556
rect 4465 3536 4469 3556
rect 4485 3536 4489 3556
rect 4505 3536 4509 3556
rect 4525 3536 4529 3556
rect 4545 3536 4549 3556
rect 4565 3536 4569 3556
rect 4465 3524 4478 3536
rect 4505 3524 4518 3536
rect 4545 3524 4558 3536
rect 4585 3533 4589 3556
rect 4605 3533 4609 3556
rect 4651 3551 4655 3556
rect 4362 3483 4371 3491
rect 4342 3464 4345 3476
rect 4335 3424 4339 3430
rect 4347 3424 4351 3464
rect 4367 3424 4371 3483
rect 4381 3424 4385 3506
rect 4401 3464 4405 3507
rect 4465 3464 4469 3524
rect 4485 3464 4489 3524
rect 4505 3464 4509 3524
rect 4525 3464 4529 3524
rect 4545 3464 4549 3524
rect 4565 3464 4569 3524
rect 4585 3521 4594 3533
rect 4606 3521 4609 3533
rect 4585 3464 4589 3521
rect 4605 3464 4609 3521
rect 4642 3544 4655 3551
rect 4642 3499 4646 3544
rect 4671 3533 4675 3556
rect 4666 3521 4675 3533
rect 4642 3476 4646 3487
rect 4642 3468 4660 3476
rect 4656 3464 4660 3468
rect 4664 3464 4668 3521
rect 4691 3479 4695 3556
rect 4686 3467 4693 3479
rect 4686 3424 4690 3467
rect 45 3380 49 3384
rect 65 3380 69 3384
rect 115 3380 119 3384
rect 135 3380 139 3384
rect 149 3380 153 3384
rect 169 3380 173 3384
rect 181 3380 185 3384
rect 201 3380 205 3384
rect 247 3380 251 3384
rect 255 3380 259 3384
rect 275 3380 279 3384
rect 283 3380 287 3384
rect 305 3380 309 3384
rect 365 3380 369 3384
rect 425 3380 429 3384
rect 445 3380 449 3384
rect 510 3380 514 3384
rect 532 3380 536 3384
rect 540 3380 544 3384
rect 610 3380 614 3384
rect 632 3380 636 3384
rect 640 3380 644 3384
rect 691 3380 695 3384
rect 711 3380 715 3384
rect 771 3380 775 3384
rect 781 3380 785 3384
rect 811 3380 815 3384
rect 821 3380 825 3384
rect 891 3380 895 3384
rect 965 3380 969 3384
rect 985 3380 989 3384
rect 1005 3380 1009 3384
rect 1051 3380 1055 3384
rect 1071 3380 1075 3384
rect 1091 3380 1095 3384
rect 1151 3380 1155 3384
rect 1159 3380 1163 3384
rect 1231 3380 1235 3384
rect 1251 3380 1255 3384
rect 1311 3380 1315 3384
rect 1331 3380 1335 3384
rect 1396 3380 1400 3384
rect 1404 3380 1408 3384
rect 1426 3380 1430 3384
rect 1495 3380 1499 3384
rect 1515 3380 1519 3384
rect 1529 3380 1533 3384
rect 1549 3380 1553 3384
rect 1561 3380 1565 3384
rect 1581 3380 1585 3384
rect 1627 3380 1631 3384
rect 1635 3380 1639 3384
rect 1655 3380 1659 3384
rect 1663 3380 1667 3384
rect 1685 3380 1689 3384
rect 1745 3380 1749 3384
rect 1765 3380 1769 3384
rect 1816 3380 1820 3384
rect 1824 3380 1828 3384
rect 1846 3380 1850 3384
rect 1911 3380 1915 3384
rect 1985 3380 1989 3384
rect 2005 3380 2009 3384
rect 2061 3380 2065 3384
rect 2083 3380 2087 3384
rect 2105 3380 2109 3384
rect 2151 3380 2155 3384
rect 2171 3380 2175 3384
rect 2231 3380 2235 3384
rect 2251 3380 2255 3384
rect 2271 3380 2275 3384
rect 2331 3380 2335 3384
rect 2391 3380 2395 3384
rect 2451 3380 2455 3384
rect 2473 3380 2477 3384
rect 2481 3380 2485 3384
rect 2501 3380 2505 3384
rect 2509 3380 2513 3384
rect 2555 3380 2559 3384
rect 2575 3380 2579 3384
rect 2587 3380 2591 3384
rect 2607 3380 2611 3384
rect 2621 3380 2625 3384
rect 2641 3380 2645 3384
rect 2696 3380 2700 3384
rect 2704 3380 2708 3384
rect 2726 3380 2730 3384
rect 2791 3380 2795 3384
rect 2813 3380 2817 3384
rect 2871 3380 2875 3384
rect 2891 3380 2895 3384
rect 2951 3380 2955 3384
rect 2973 3380 2977 3384
rect 2981 3380 2985 3384
rect 3001 3380 3005 3384
rect 3009 3380 3013 3384
rect 3055 3380 3059 3384
rect 3075 3380 3079 3384
rect 3087 3380 3091 3384
rect 3107 3380 3111 3384
rect 3121 3380 3125 3384
rect 3141 3380 3145 3384
rect 3210 3380 3214 3384
rect 3232 3380 3236 3384
rect 3240 3380 3244 3384
rect 3305 3380 3309 3384
rect 3351 3380 3355 3384
rect 3359 3380 3363 3384
rect 3431 3380 3435 3384
rect 3517 3380 3521 3384
rect 3525 3380 3529 3384
rect 3571 3380 3575 3384
rect 3591 3380 3595 3384
rect 3611 3380 3615 3384
rect 3671 3380 3675 3384
rect 3681 3380 3685 3384
rect 3701 3380 3705 3384
rect 3785 3380 3789 3384
rect 3805 3380 3809 3384
rect 3825 3380 3829 3384
rect 3845 3380 3849 3384
rect 3905 3380 3909 3384
rect 3925 3380 3929 3384
rect 3971 3380 3975 3384
rect 3993 3380 3997 3384
rect 4001 3380 4005 3384
rect 4021 3380 4025 3384
rect 4029 3380 4033 3384
rect 4075 3380 4079 3384
rect 4095 3380 4099 3384
rect 4107 3380 4111 3384
rect 4127 3380 4131 3384
rect 4141 3380 4145 3384
rect 4161 3380 4165 3384
rect 4211 3380 4215 3384
rect 4233 3380 4237 3384
rect 4241 3380 4245 3384
rect 4261 3380 4265 3384
rect 4269 3380 4273 3384
rect 4315 3380 4319 3384
rect 4335 3380 4339 3384
rect 4347 3380 4351 3384
rect 4367 3380 4371 3384
rect 4381 3380 4385 3384
rect 4401 3380 4405 3384
rect 4465 3380 4469 3384
rect 4485 3380 4489 3384
rect 4505 3380 4509 3384
rect 4525 3380 4529 3384
rect 4545 3380 4549 3384
rect 4565 3380 4569 3384
rect 4585 3380 4589 3384
rect 4605 3380 4609 3384
rect 4656 3380 4660 3384
rect 4664 3380 4668 3384
rect 4686 3380 4690 3384
rect 35 3356 39 3360
rect 55 3356 59 3360
rect 69 3356 73 3360
rect 89 3356 93 3360
rect 101 3356 105 3360
rect 121 3356 125 3360
rect 167 3356 171 3360
rect 175 3356 179 3360
rect 195 3356 199 3360
rect 203 3356 207 3360
rect 225 3356 229 3360
rect 285 3356 289 3360
rect 305 3356 309 3360
rect 325 3356 329 3360
rect 345 3356 349 3360
rect 405 3356 409 3360
rect 425 3356 429 3360
rect 471 3356 475 3360
rect 493 3356 497 3360
rect 501 3356 505 3360
rect 521 3356 525 3360
rect 529 3356 533 3360
rect 575 3356 579 3360
rect 595 3356 599 3360
rect 607 3356 611 3360
rect 627 3356 631 3360
rect 641 3356 645 3360
rect 661 3356 665 3360
rect 730 3356 734 3360
rect 752 3356 756 3360
rect 760 3356 764 3360
rect 825 3356 829 3360
rect 845 3356 849 3360
rect 865 3356 869 3360
rect 885 3356 889 3360
rect 931 3356 935 3360
rect 951 3356 955 3360
rect 1025 3356 1029 3360
rect 1045 3356 1049 3360
rect 1065 3356 1069 3360
rect 1121 3356 1125 3360
rect 1143 3356 1147 3360
rect 1165 3356 1169 3360
rect 1211 3356 1215 3360
rect 1231 3356 1235 3360
rect 1251 3356 1255 3360
rect 1316 3356 1320 3360
rect 1324 3356 1328 3360
rect 1346 3356 1350 3360
rect 1411 3356 1415 3360
rect 1431 3356 1435 3360
rect 1515 3356 1519 3360
rect 1535 3356 1539 3360
rect 1545 3356 1549 3360
rect 1605 3356 1609 3360
rect 1625 3356 1629 3360
rect 1676 3356 1680 3360
rect 1684 3356 1688 3360
rect 1706 3356 1710 3360
rect 1790 3356 1794 3360
rect 1812 3356 1816 3360
rect 1820 3356 1824 3360
rect 1871 3356 1875 3360
rect 1891 3356 1895 3360
rect 1956 3356 1960 3360
rect 1964 3356 1968 3360
rect 1986 3356 1990 3360
rect 2070 3356 2074 3360
rect 2092 3356 2096 3360
rect 2100 3356 2104 3360
rect 2151 3356 2155 3360
rect 2216 3356 2220 3360
rect 2224 3356 2228 3360
rect 2246 3356 2250 3360
rect 2325 3356 2329 3360
rect 2371 3356 2375 3360
rect 2391 3356 2395 3360
rect 2451 3356 2455 3360
rect 2473 3356 2477 3360
rect 2481 3356 2485 3360
rect 2501 3356 2505 3360
rect 2509 3356 2513 3360
rect 2555 3356 2559 3360
rect 2575 3356 2579 3360
rect 2587 3356 2591 3360
rect 2607 3356 2611 3360
rect 2621 3356 2625 3360
rect 2641 3356 2645 3360
rect 2691 3356 2695 3360
rect 2713 3356 2717 3360
rect 2771 3356 2775 3360
rect 2793 3356 2797 3360
rect 2801 3356 2805 3360
rect 2821 3356 2825 3360
rect 2829 3356 2833 3360
rect 2875 3356 2879 3360
rect 2895 3356 2899 3360
rect 2907 3356 2911 3360
rect 2927 3356 2931 3360
rect 2941 3356 2945 3360
rect 2961 3356 2965 3360
rect 3030 3356 3034 3360
rect 3052 3356 3056 3360
rect 3060 3356 3064 3360
rect 3130 3356 3134 3360
rect 3152 3356 3156 3360
rect 3160 3356 3164 3360
rect 3216 3356 3220 3360
rect 3224 3356 3228 3360
rect 3246 3356 3250 3360
rect 3330 3356 3334 3360
rect 3352 3356 3356 3360
rect 3360 3356 3364 3360
rect 3416 3356 3420 3360
rect 3424 3356 3428 3360
rect 3446 3356 3450 3360
rect 3511 3356 3515 3360
rect 3531 3356 3535 3360
rect 3591 3356 3595 3360
rect 3611 3356 3615 3360
rect 3671 3356 3675 3360
rect 3691 3356 3695 3360
rect 3751 3356 3755 3360
rect 3771 3356 3775 3360
rect 3831 3356 3835 3360
rect 3853 3356 3857 3360
rect 3925 3356 3929 3360
rect 3945 3356 3949 3360
rect 4017 3356 4021 3360
rect 4025 3356 4029 3360
rect 4071 3356 4075 3360
rect 4093 3356 4097 3360
rect 4165 3356 4169 3360
rect 4230 3356 4234 3360
rect 4252 3356 4256 3360
rect 4260 3356 4264 3360
rect 4325 3356 4329 3360
rect 4376 3356 4380 3360
rect 4384 3356 4388 3360
rect 4406 3356 4410 3360
rect 4485 3356 4489 3360
rect 4505 3356 4509 3360
rect 4555 3356 4559 3360
rect 4575 3356 4579 3360
rect 4589 3356 4593 3360
rect 4609 3356 4613 3360
rect 4621 3356 4625 3360
rect 4641 3356 4645 3360
rect 4687 3356 4691 3360
rect 4695 3356 4699 3360
rect 4715 3356 4719 3360
rect 4723 3356 4727 3360
rect 4745 3356 4749 3360
rect 35 3233 39 3276
rect 55 3234 59 3316
rect 69 3257 73 3316
rect 89 3276 93 3316
rect 101 3310 105 3316
rect 95 3264 98 3276
rect 69 3249 78 3257
rect 35 3184 39 3221
rect 55 3164 59 3222
rect 74 3220 78 3249
rect 94 3200 98 3264
rect 65 3196 98 3200
rect 65 3164 69 3196
rect 103 3188 107 3298
rect 121 3290 125 3316
rect 167 3312 171 3316
rect 135 3310 171 3312
rect 147 3308 171 3310
rect 89 3176 91 3188
rect 87 3164 91 3176
rect 97 3176 99 3188
rect 97 3164 101 3176
rect 119 3164 123 3278
rect 135 3172 139 3298
rect 175 3284 179 3316
rect 195 3296 199 3336
rect 203 3313 207 3336
rect 203 3306 211 3313
rect 173 3189 179 3284
rect 207 3277 211 3306
rect 203 3271 211 3277
rect 203 3225 207 3271
rect 225 3264 229 3276
rect 227 3252 229 3264
rect 285 3253 289 3276
rect 173 3185 197 3189
rect 159 3180 177 3181
rect 147 3176 177 3180
rect 135 3168 169 3172
rect 165 3164 169 3168
rect 173 3164 177 3176
rect 193 3164 197 3185
rect 203 3164 207 3213
rect 225 3184 229 3252
rect 286 3241 289 3253
rect 280 3193 286 3241
rect 305 3219 309 3276
rect 325 3254 329 3276
rect 345 3254 349 3276
rect 325 3248 338 3254
rect 345 3253 365 3254
rect 345 3248 353 3253
rect 334 3219 338 3248
rect 307 3207 309 3219
rect 305 3205 309 3207
rect 305 3198 318 3205
rect 280 3189 310 3193
rect 306 3184 310 3189
rect 314 3184 318 3198
rect 334 3184 338 3207
rect 353 3199 359 3241
rect 405 3239 409 3316
rect 406 3227 409 3239
rect 403 3211 409 3227
rect 425 3239 429 3316
rect 493 3313 497 3336
rect 489 3306 497 3313
rect 489 3277 493 3306
rect 501 3296 505 3336
rect 521 3284 525 3316
rect 529 3312 533 3316
rect 529 3310 565 3312
rect 529 3308 553 3310
rect 471 3264 475 3276
rect 489 3271 497 3277
rect 471 3252 473 3264
rect 425 3227 434 3239
rect 425 3211 431 3227
rect 403 3204 417 3211
rect 342 3192 359 3199
rect 342 3184 346 3192
rect 413 3184 417 3204
rect 423 3204 431 3211
rect 423 3184 427 3204
rect 471 3184 475 3252
rect 493 3225 497 3271
rect 493 3164 497 3213
rect 521 3189 527 3284
rect 503 3185 527 3189
rect 503 3164 507 3185
rect 523 3180 541 3181
rect 523 3176 553 3180
rect 523 3164 527 3176
rect 561 3172 565 3298
rect 575 3290 579 3316
rect 595 3310 599 3316
rect 531 3168 565 3172
rect 531 3164 535 3168
rect 577 3164 581 3278
rect 593 3188 597 3298
rect 607 3276 611 3316
rect 602 3264 605 3276
rect 602 3200 606 3264
rect 627 3257 631 3316
rect 622 3249 631 3257
rect 622 3220 626 3249
rect 641 3234 645 3316
rect 661 3233 665 3276
rect 730 3273 734 3316
rect 727 3261 734 3273
rect 602 3196 635 3200
rect 601 3176 603 3188
rect 599 3164 603 3176
rect 609 3176 611 3188
rect 609 3164 613 3176
rect 631 3164 635 3196
rect 641 3164 645 3222
rect 661 3184 665 3221
rect 725 3184 729 3261
rect 752 3219 756 3276
rect 760 3272 764 3276
rect 760 3264 778 3272
rect 774 3253 778 3264
rect 825 3253 829 3276
rect 826 3241 829 3253
rect 745 3207 754 3219
rect 745 3184 749 3207
rect 774 3196 778 3241
rect 765 3189 778 3196
rect 820 3193 826 3241
rect 845 3219 849 3276
rect 865 3254 869 3276
rect 885 3254 889 3276
rect 865 3248 878 3254
rect 885 3253 905 3254
rect 885 3248 893 3253
rect 874 3219 878 3248
rect 847 3207 849 3219
rect 845 3205 849 3207
rect 845 3198 858 3205
rect 820 3189 850 3193
rect 765 3184 769 3189
rect 846 3184 850 3189
rect 854 3184 858 3198
rect 874 3184 878 3207
rect 893 3199 899 3241
rect 931 3239 935 3316
rect 926 3227 935 3239
rect 929 3211 935 3227
rect 951 3239 955 3316
rect 1025 3273 1029 3316
rect 1045 3304 1049 3316
rect 1065 3308 1069 3316
rect 1065 3304 1080 3308
rect 1045 3300 1060 3304
rect 1054 3293 1060 3300
rect 1025 3261 1033 3273
rect 1045 3261 1052 3273
rect 951 3227 954 3239
rect 951 3211 957 3227
rect 929 3204 937 3211
rect 882 3192 899 3199
rect 882 3184 886 3192
rect 933 3184 937 3204
rect 943 3204 957 3211
rect 1048 3204 1052 3261
rect 1056 3204 1060 3281
rect 1074 3273 1080 3304
rect 1064 3261 1074 3273
rect 1064 3204 1068 3261
rect 943 3184 947 3204
rect 1121 3202 1125 3276
rect 1143 3239 1147 3316
rect 1165 3253 1169 3316
rect 1211 3308 1215 3316
rect 1200 3304 1215 3308
rect 1231 3304 1235 3316
rect 1200 3273 1206 3304
rect 1220 3300 1235 3304
rect 1220 3293 1226 3300
rect 1206 3261 1216 3273
rect 1165 3241 1174 3253
rect 1146 3227 1159 3239
rect 1121 3190 1133 3202
rect 1135 3184 1139 3190
rect 1155 3184 1159 3227
rect 1165 3184 1169 3241
rect 1212 3204 1216 3261
rect 1220 3204 1224 3281
rect 1251 3273 1255 3316
rect 1228 3261 1235 3273
rect 1247 3261 1255 3273
rect 1316 3272 1320 3276
rect 1302 3264 1320 3272
rect 1228 3204 1232 3261
rect 1302 3253 1306 3264
rect 1302 3196 1306 3241
rect 1324 3219 1328 3276
rect 1346 3273 1350 3316
rect 1346 3261 1353 3273
rect 1326 3207 1335 3219
rect 1302 3189 1315 3196
rect 1311 3184 1315 3189
rect 1331 3184 1335 3207
rect 1351 3184 1355 3261
rect 1411 3239 1415 3316
rect 1406 3227 1415 3239
rect 1409 3211 1415 3227
rect 1431 3239 1435 3316
rect 1515 3271 1519 3276
rect 1535 3253 1539 3276
rect 1545 3272 1549 3276
rect 1545 3267 1558 3272
rect 1431 3227 1434 3239
rect 1431 3211 1437 3227
rect 1409 3204 1417 3211
rect 1413 3184 1417 3204
rect 1423 3204 1437 3211
rect 1423 3184 1427 3204
rect 1505 3192 1515 3204
rect 1505 3184 1509 3192
rect 1535 3177 1539 3241
rect 1525 3171 1539 3177
rect 1554 3233 1558 3267
rect 1605 3239 1609 3316
rect 1606 3227 1609 3239
rect 1554 3176 1558 3221
rect 1603 3211 1609 3227
rect 1625 3239 1629 3316
rect 1676 3272 1680 3276
rect 1662 3264 1680 3272
rect 1662 3253 1666 3264
rect 1625 3227 1634 3239
rect 1625 3211 1631 3227
rect 1603 3204 1617 3211
rect 1613 3184 1617 3204
rect 1623 3204 1631 3211
rect 1623 3184 1627 3204
rect 1662 3196 1666 3241
rect 1684 3219 1688 3276
rect 1706 3273 1710 3316
rect 1790 3273 1794 3316
rect 1706 3261 1713 3273
rect 1787 3261 1794 3273
rect 1686 3207 1695 3219
rect 1662 3189 1675 3196
rect 1671 3184 1675 3189
rect 1691 3184 1695 3207
rect 1711 3184 1715 3261
rect 1785 3184 1789 3261
rect 1812 3219 1816 3276
rect 1820 3272 1824 3276
rect 1820 3264 1838 3272
rect 1834 3253 1838 3264
rect 1805 3207 1814 3219
rect 1805 3184 1809 3207
rect 1834 3196 1838 3241
rect 1871 3239 1875 3316
rect 1866 3227 1875 3239
rect 1869 3211 1875 3227
rect 1891 3239 1895 3316
rect 1956 3272 1960 3276
rect 1942 3264 1960 3272
rect 1942 3253 1946 3264
rect 1891 3227 1894 3239
rect 1891 3211 1897 3227
rect 1869 3204 1877 3211
rect 1825 3189 1838 3196
rect 1825 3184 1829 3189
rect 1873 3184 1877 3204
rect 1883 3204 1897 3211
rect 1883 3184 1887 3204
rect 1942 3196 1946 3241
rect 1964 3219 1968 3276
rect 1986 3273 1990 3316
rect 2070 3273 2074 3316
rect 1986 3261 1993 3273
rect 2067 3261 2074 3273
rect 1966 3207 1975 3219
rect 1942 3189 1955 3196
rect 1951 3184 1955 3189
rect 1971 3184 1975 3207
rect 1991 3184 1995 3261
rect 2065 3184 2069 3261
rect 2092 3219 2096 3276
rect 2100 3272 2104 3276
rect 2100 3264 2118 3272
rect 2114 3253 2118 3264
rect 2085 3207 2094 3219
rect 2085 3184 2089 3207
rect 2114 3196 2118 3241
rect 2151 3233 2155 3316
rect 2216 3272 2220 3276
rect 2202 3264 2220 3272
rect 2202 3253 2206 3264
rect 2146 3221 2155 3233
rect 2105 3189 2118 3196
rect 2105 3184 2109 3189
rect 1545 3171 1558 3176
rect 1525 3164 1529 3171
rect 1545 3164 1549 3171
rect 2151 3164 2155 3221
rect 2202 3196 2206 3241
rect 2224 3219 2228 3276
rect 2246 3273 2250 3316
rect 2246 3261 2253 3273
rect 2226 3207 2235 3219
rect 2202 3189 2215 3196
rect 2211 3184 2215 3189
rect 2231 3184 2235 3207
rect 2251 3184 2255 3261
rect 2325 3233 2329 3316
rect 2371 3239 2375 3316
rect 2325 3221 2334 3233
rect 2366 3227 2375 3239
rect 2325 3164 2329 3221
rect 2369 3211 2375 3227
rect 2391 3239 2395 3316
rect 2473 3313 2477 3336
rect 2469 3306 2477 3313
rect 2469 3277 2473 3306
rect 2481 3296 2485 3336
rect 2501 3284 2505 3316
rect 2509 3312 2513 3316
rect 2509 3310 2545 3312
rect 2509 3308 2533 3310
rect 2451 3264 2455 3276
rect 2469 3271 2477 3277
rect 2451 3252 2453 3264
rect 2391 3227 2394 3239
rect 2391 3211 2397 3227
rect 2369 3204 2377 3211
rect 2373 3184 2377 3204
rect 2383 3204 2397 3211
rect 2383 3184 2387 3204
rect 2451 3184 2455 3252
rect 2473 3225 2477 3271
rect 2473 3164 2477 3213
rect 2501 3189 2507 3284
rect 2483 3185 2507 3189
rect 2483 3164 2487 3185
rect 2503 3180 2521 3181
rect 2503 3176 2533 3180
rect 2503 3164 2507 3176
rect 2541 3172 2545 3298
rect 2555 3290 2559 3316
rect 2575 3310 2579 3316
rect 2511 3168 2545 3172
rect 2511 3164 2515 3168
rect 2557 3164 2561 3278
rect 2573 3188 2577 3298
rect 2587 3276 2591 3316
rect 2582 3264 2585 3276
rect 2582 3200 2586 3264
rect 2607 3257 2611 3316
rect 2602 3249 2611 3257
rect 2602 3220 2606 3249
rect 2621 3234 2625 3316
rect 2641 3233 2645 3276
rect 2691 3253 2695 3316
rect 2793 3313 2797 3336
rect 2789 3306 2797 3313
rect 2789 3277 2793 3306
rect 2801 3296 2805 3336
rect 2821 3284 2825 3316
rect 2829 3312 2833 3316
rect 2829 3310 2865 3312
rect 2829 3308 2853 3310
rect 2713 3270 2717 3276
rect 2715 3258 2717 3270
rect 2771 3264 2775 3276
rect 2789 3271 2797 3277
rect 2686 3241 2695 3253
rect 2582 3196 2615 3200
rect 2581 3176 2583 3188
rect 2579 3164 2583 3176
rect 2589 3176 2591 3188
rect 2589 3164 2593 3176
rect 2611 3164 2615 3196
rect 2621 3164 2625 3222
rect 2641 3184 2645 3221
rect 2691 3164 2695 3241
rect 2771 3252 2773 3264
rect 2715 3190 2717 3202
rect 2713 3184 2717 3190
rect 2771 3184 2775 3252
rect 2793 3225 2797 3271
rect 2793 3164 2797 3213
rect 2821 3189 2827 3284
rect 2803 3185 2827 3189
rect 2803 3164 2807 3185
rect 2823 3180 2841 3181
rect 2823 3176 2853 3180
rect 2823 3164 2827 3176
rect 2861 3172 2865 3298
rect 2875 3290 2879 3316
rect 2895 3310 2899 3316
rect 2831 3168 2865 3172
rect 2831 3164 2835 3168
rect 2877 3164 2881 3278
rect 2893 3188 2897 3298
rect 2907 3276 2911 3316
rect 2902 3264 2905 3276
rect 2902 3200 2906 3264
rect 2927 3257 2931 3316
rect 2922 3249 2931 3257
rect 2922 3220 2926 3249
rect 2941 3234 2945 3316
rect 2961 3233 2965 3276
rect 3030 3273 3034 3316
rect 3027 3261 3034 3273
rect 2902 3196 2935 3200
rect 2901 3176 2903 3188
rect 2899 3164 2903 3176
rect 2909 3176 2911 3188
rect 2909 3164 2913 3176
rect 2931 3164 2935 3196
rect 2941 3164 2945 3222
rect 2961 3184 2965 3221
rect 3025 3184 3029 3261
rect 3052 3219 3056 3276
rect 3060 3272 3064 3276
rect 3130 3273 3134 3316
rect 3060 3264 3078 3272
rect 3074 3253 3078 3264
rect 3127 3261 3134 3273
rect 3045 3207 3054 3219
rect 3045 3184 3049 3207
rect 3074 3196 3078 3241
rect 3065 3189 3078 3196
rect 3065 3184 3069 3189
rect 3125 3184 3129 3261
rect 3152 3219 3156 3276
rect 3160 3272 3164 3276
rect 3216 3272 3220 3276
rect 3160 3264 3178 3272
rect 3174 3253 3178 3264
rect 3202 3264 3220 3272
rect 3202 3253 3206 3264
rect 3145 3207 3154 3219
rect 3145 3184 3149 3207
rect 3174 3196 3178 3241
rect 3165 3189 3178 3196
rect 3202 3196 3206 3241
rect 3224 3219 3228 3276
rect 3246 3273 3250 3316
rect 3330 3273 3334 3316
rect 3246 3261 3253 3273
rect 3327 3261 3334 3273
rect 3226 3207 3235 3219
rect 3202 3189 3215 3196
rect 3165 3184 3169 3189
rect 3211 3184 3215 3189
rect 3231 3184 3235 3207
rect 3251 3184 3255 3261
rect 3325 3184 3329 3261
rect 3352 3219 3356 3276
rect 3360 3272 3364 3276
rect 3416 3272 3420 3276
rect 3360 3264 3378 3272
rect 3374 3253 3378 3264
rect 3402 3264 3420 3272
rect 3402 3253 3406 3264
rect 3345 3207 3354 3219
rect 3345 3184 3349 3207
rect 3374 3196 3378 3241
rect 3365 3189 3378 3196
rect 3402 3196 3406 3241
rect 3424 3219 3428 3276
rect 3446 3273 3450 3316
rect 3446 3261 3453 3273
rect 3426 3207 3435 3219
rect 3402 3189 3415 3196
rect 3365 3184 3369 3189
rect 3411 3184 3415 3189
rect 3431 3184 3435 3207
rect 3451 3184 3455 3261
rect 3511 3239 3515 3316
rect 3506 3227 3515 3239
rect 3509 3211 3515 3227
rect 3531 3239 3535 3316
rect 3591 3239 3595 3316
rect 3531 3227 3534 3239
rect 3586 3227 3595 3239
rect 3531 3211 3537 3227
rect 3509 3204 3517 3211
rect 3513 3184 3517 3204
rect 3523 3204 3537 3211
rect 3589 3211 3595 3227
rect 3611 3239 3615 3316
rect 3671 3239 3675 3316
rect 3611 3227 3614 3239
rect 3666 3227 3675 3239
rect 3611 3211 3617 3227
rect 3589 3204 3597 3211
rect 3523 3184 3527 3204
rect 3593 3184 3597 3204
rect 3603 3204 3617 3211
rect 3669 3211 3675 3227
rect 3691 3239 3695 3316
rect 3751 3239 3755 3316
rect 3691 3227 3694 3239
rect 3746 3227 3755 3239
rect 3691 3211 3697 3227
rect 3669 3204 3677 3211
rect 3603 3184 3607 3204
rect 3673 3184 3677 3204
rect 3683 3204 3697 3211
rect 3749 3211 3755 3227
rect 3771 3239 3775 3316
rect 3831 3253 3835 3316
rect 3853 3270 3857 3276
rect 3855 3258 3857 3270
rect 3826 3241 3835 3253
rect 3771 3227 3774 3239
rect 3771 3211 3777 3227
rect 3749 3204 3757 3211
rect 3683 3184 3687 3204
rect 3753 3184 3757 3204
rect 3763 3204 3777 3211
rect 3763 3184 3767 3204
rect 3831 3164 3835 3241
rect 3925 3239 3929 3316
rect 3926 3227 3929 3239
rect 3923 3211 3929 3227
rect 3945 3239 3949 3316
rect 4017 3253 4021 3276
rect 4006 3241 4021 3253
rect 4025 3253 4029 3276
rect 4071 3253 4075 3316
rect 4093 3270 4097 3276
rect 4095 3258 4097 3270
rect 4025 3241 4034 3253
rect 4066 3241 4075 3253
rect 3945 3227 3954 3239
rect 3945 3211 3951 3227
rect 3923 3204 3937 3211
rect 3855 3190 3857 3202
rect 3853 3184 3857 3190
rect 3933 3184 3937 3204
rect 3943 3204 3951 3211
rect 3943 3184 3947 3204
rect 4005 3164 4009 3241
rect 4025 3164 4029 3241
rect 4071 3164 4075 3241
rect 4165 3233 4169 3316
rect 4230 3273 4234 3316
rect 4227 3261 4234 3273
rect 4165 3221 4174 3233
rect 4095 3190 4097 3202
rect 4093 3184 4097 3190
rect 4165 3164 4169 3221
rect 4225 3184 4229 3261
rect 4252 3219 4256 3276
rect 4260 3272 4264 3276
rect 4260 3264 4278 3272
rect 4274 3253 4278 3264
rect 4245 3207 4254 3219
rect 4245 3184 4249 3207
rect 4274 3196 4278 3241
rect 4265 3189 4278 3196
rect 4325 3233 4329 3316
rect 4376 3272 4380 3276
rect 4362 3264 4380 3272
rect 4362 3253 4366 3264
rect 4325 3221 4334 3233
rect 4265 3184 4269 3189
rect 4325 3164 4329 3221
rect 4362 3196 4366 3241
rect 4384 3219 4388 3276
rect 4406 3273 4410 3316
rect 4406 3261 4413 3273
rect 4386 3207 4395 3219
rect 4362 3189 4375 3196
rect 4371 3184 4375 3189
rect 4391 3184 4395 3207
rect 4411 3184 4415 3261
rect 4485 3239 4489 3316
rect 4486 3227 4489 3239
rect 4483 3211 4489 3227
rect 4505 3239 4509 3316
rect 4505 3227 4514 3239
rect 4555 3233 4559 3276
rect 4575 3234 4579 3316
rect 4589 3257 4593 3316
rect 4609 3276 4613 3316
rect 4621 3310 4625 3316
rect 4615 3264 4618 3276
rect 4589 3249 4598 3257
rect 4505 3211 4511 3227
rect 4483 3204 4497 3211
rect 4493 3184 4497 3204
rect 4503 3204 4511 3211
rect 4503 3184 4507 3204
rect 4555 3184 4559 3221
rect 4575 3164 4579 3222
rect 4594 3220 4598 3249
rect 4614 3200 4618 3264
rect 4585 3196 4618 3200
rect 4585 3164 4589 3196
rect 4623 3188 4627 3298
rect 4641 3290 4645 3316
rect 4687 3312 4691 3316
rect 4655 3310 4691 3312
rect 4667 3308 4691 3310
rect 4609 3176 4611 3188
rect 4607 3164 4611 3176
rect 4617 3176 4619 3188
rect 4617 3164 4621 3176
rect 4639 3164 4643 3278
rect 4655 3172 4659 3298
rect 4695 3284 4699 3316
rect 4715 3296 4719 3336
rect 4723 3313 4727 3336
rect 4723 3306 4731 3313
rect 4693 3189 4699 3284
rect 4727 3277 4731 3306
rect 4723 3271 4731 3277
rect 4723 3225 4727 3271
rect 4745 3264 4749 3276
rect 4747 3252 4749 3264
rect 4693 3185 4717 3189
rect 4679 3180 4697 3181
rect 4667 3176 4697 3180
rect 4655 3168 4689 3172
rect 4685 3164 4689 3168
rect 4693 3164 4697 3176
rect 4713 3164 4717 3185
rect 4723 3164 4727 3213
rect 4745 3184 4749 3252
rect 35 3140 39 3144
rect 55 3140 59 3144
rect 65 3140 69 3144
rect 87 3140 91 3144
rect 97 3140 101 3144
rect 119 3140 123 3144
rect 165 3140 169 3144
rect 173 3140 177 3144
rect 193 3140 197 3144
rect 203 3140 207 3144
rect 225 3140 229 3144
rect 306 3140 310 3144
rect 314 3140 318 3144
rect 334 3140 338 3144
rect 342 3140 346 3144
rect 413 3140 417 3144
rect 423 3140 427 3144
rect 471 3140 475 3144
rect 493 3140 497 3144
rect 503 3140 507 3144
rect 523 3140 527 3144
rect 531 3140 535 3144
rect 577 3140 581 3144
rect 599 3140 603 3144
rect 609 3140 613 3144
rect 631 3140 635 3144
rect 641 3140 645 3144
rect 661 3140 665 3144
rect 725 3140 729 3144
rect 745 3140 749 3144
rect 765 3140 769 3144
rect 846 3140 850 3144
rect 854 3140 858 3144
rect 874 3140 878 3144
rect 882 3140 886 3144
rect 933 3140 937 3144
rect 943 3140 947 3144
rect 1048 3140 1052 3144
rect 1056 3140 1060 3144
rect 1064 3140 1068 3144
rect 1135 3140 1139 3144
rect 1155 3140 1159 3144
rect 1165 3140 1169 3144
rect 1212 3140 1216 3144
rect 1220 3140 1224 3144
rect 1228 3140 1232 3144
rect 1311 3140 1315 3144
rect 1331 3140 1335 3144
rect 1351 3140 1355 3144
rect 1413 3140 1417 3144
rect 1423 3140 1427 3144
rect 1505 3140 1509 3144
rect 1525 3140 1529 3144
rect 1545 3140 1549 3144
rect 1613 3140 1617 3144
rect 1623 3140 1627 3144
rect 1671 3140 1675 3144
rect 1691 3140 1695 3144
rect 1711 3140 1715 3144
rect 1785 3140 1789 3144
rect 1805 3140 1809 3144
rect 1825 3140 1829 3144
rect 1873 3140 1877 3144
rect 1883 3140 1887 3144
rect 1951 3140 1955 3144
rect 1971 3140 1975 3144
rect 1991 3140 1995 3144
rect 2065 3140 2069 3144
rect 2085 3140 2089 3144
rect 2105 3140 2109 3144
rect 2151 3140 2155 3144
rect 2211 3140 2215 3144
rect 2231 3140 2235 3144
rect 2251 3140 2255 3144
rect 2325 3140 2329 3144
rect 2373 3140 2377 3144
rect 2383 3140 2387 3144
rect 2451 3140 2455 3144
rect 2473 3140 2477 3144
rect 2483 3140 2487 3144
rect 2503 3140 2507 3144
rect 2511 3140 2515 3144
rect 2557 3140 2561 3144
rect 2579 3140 2583 3144
rect 2589 3140 2593 3144
rect 2611 3140 2615 3144
rect 2621 3140 2625 3144
rect 2641 3140 2645 3144
rect 2691 3140 2695 3144
rect 2713 3140 2717 3144
rect 2771 3140 2775 3144
rect 2793 3140 2797 3144
rect 2803 3140 2807 3144
rect 2823 3140 2827 3144
rect 2831 3140 2835 3144
rect 2877 3140 2881 3144
rect 2899 3140 2903 3144
rect 2909 3140 2913 3144
rect 2931 3140 2935 3144
rect 2941 3140 2945 3144
rect 2961 3140 2965 3144
rect 3025 3140 3029 3144
rect 3045 3140 3049 3144
rect 3065 3140 3069 3144
rect 3125 3140 3129 3144
rect 3145 3140 3149 3144
rect 3165 3140 3169 3144
rect 3211 3140 3215 3144
rect 3231 3140 3235 3144
rect 3251 3140 3255 3144
rect 3325 3140 3329 3144
rect 3345 3140 3349 3144
rect 3365 3140 3369 3144
rect 3411 3140 3415 3144
rect 3431 3140 3435 3144
rect 3451 3140 3455 3144
rect 3513 3140 3517 3144
rect 3523 3140 3527 3144
rect 3593 3140 3597 3144
rect 3603 3140 3607 3144
rect 3673 3140 3677 3144
rect 3683 3140 3687 3144
rect 3753 3140 3757 3144
rect 3763 3140 3767 3144
rect 3831 3140 3835 3144
rect 3853 3140 3857 3144
rect 3933 3140 3937 3144
rect 3943 3140 3947 3144
rect 4005 3140 4009 3144
rect 4025 3140 4029 3144
rect 4071 3140 4075 3144
rect 4093 3140 4097 3144
rect 4165 3140 4169 3144
rect 4225 3140 4229 3144
rect 4245 3140 4249 3144
rect 4265 3140 4269 3144
rect 4325 3140 4329 3144
rect 4371 3140 4375 3144
rect 4391 3140 4395 3144
rect 4411 3140 4415 3144
rect 4493 3140 4497 3144
rect 4503 3140 4507 3144
rect 4555 3140 4559 3144
rect 4575 3140 4579 3144
rect 4585 3140 4589 3144
rect 4607 3140 4611 3144
rect 4617 3140 4621 3144
rect 4639 3140 4643 3144
rect 4685 3140 4689 3144
rect 4693 3140 4697 3144
rect 4713 3140 4717 3144
rect 4723 3140 4727 3144
rect 4745 3140 4749 3144
rect 66 3116 70 3120
rect 74 3116 78 3120
rect 94 3116 98 3120
rect 102 3116 106 3120
rect 175 3116 179 3120
rect 195 3116 199 3120
rect 205 3116 209 3120
rect 251 3116 255 3120
rect 273 3116 277 3120
rect 283 3116 287 3120
rect 303 3116 307 3120
rect 311 3116 315 3120
rect 357 3116 361 3120
rect 379 3116 383 3120
rect 389 3116 393 3120
rect 411 3116 415 3120
rect 421 3116 425 3120
rect 441 3116 445 3120
rect 491 3116 495 3120
rect 511 3116 515 3120
rect 531 3116 535 3120
rect 593 3116 597 3120
rect 603 3116 607 3120
rect 693 3116 697 3120
rect 703 3116 707 3120
rect 765 3116 769 3120
rect 785 3116 789 3120
rect 833 3116 837 3120
rect 843 3116 847 3120
rect 925 3116 929 3120
rect 945 3116 949 3120
rect 965 3116 969 3120
rect 1025 3116 1029 3120
rect 1045 3116 1049 3120
rect 1065 3116 1069 3120
rect 1125 3116 1129 3120
rect 1145 3116 1149 3120
rect 1205 3116 1209 3120
rect 1225 3116 1229 3120
rect 1245 3116 1249 3120
rect 1293 3116 1297 3120
rect 1303 3116 1307 3120
rect 1385 3116 1389 3120
rect 1433 3116 1437 3120
rect 1443 3116 1447 3120
rect 1513 3116 1517 3120
rect 1523 3116 1527 3120
rect 1591 3116 1595 3120
rect 1613 3116 1617 3120
rect 1671 3116 1675 3120
rect 1691 3116 1695 3120
rect 1711 3116 1715 3120
rect 1771 3116 1775 3120
rect 1791 3116 1795 3120
rect 1811 3116 1815 3120
rect 1871 3116 1875 3120
rect 1891 3116 1895 3120
rect 1954 3116 1958 3120
rect 1962 3116 1966 3120
rect 1984 3116 1988 3120
rect 2051 3116 2055 3120
rect 2111 3116 2115 3120
rect 2131 3116 2135 3120
rect 2151 3116 2155 3120
rect 2211 3116 2215 3120
rect 2231 3116 2235 3120
rect 2313 3116 2317 3120
rect 2323 3116 2327 3120
rect 2371 3116 2375 3120
rect 2391 3116 2395 3120
rect 2411 3116 2415 3120
rect 2471 3116 2475 3120
rect 2531 3116 2535 3120
rect 2551 3116 2555 3120
rect 2571 3116 2575 3120
rect 2631 3116 2635 3120
rect 2653 3116 2657 3120
rect 2713 3116 2717 3120
rect 2723 3116 2727 3120
rect 2795 3116 2799 3120
rect 2815 3116 2819 3120
rect 2825 3116 2829 3120
rect 2847 3116 2851 3120
rect 2857 3116 2861 3120
rect 2879 3116 2883 3120
rect 2925 3116 2929 3120
rect 2933 3116 2937 3120
rect 2953 3116 2957 3120
rect 2963 3116 2967 3120
rect 2985 3116 2989 3120
rect 3045 3116 3049 3120
rect 3065 3116 3069 3120
rect 3132 3116 3136 3120
rect 3154 3116 3158 3120
rect 3162 3116 3166 3120
rect 3211 3116 3215 3120
rect 3231 3116 3235 3120
rect 3295 3116 3299 3120
rect 3315 3116 3319 3120
rect 3325 3116 3329 3120
rect 3347 3116 3351 3120
rect 3357 3116 3361 3120
rect 3379 3116 3383 3120
rect 3425 3116 3429 3120
rect 3433 3116 3437 3120
rect 3453 3116 3457 3120
rect 3463 3116 3467 3120
rect 3485 3116 3489 3120
rect 3535 3116 3539 3120
rect 3555 3116 3559 3120
rect 3565 3116 3569 3120
rect 3587 3116 3591 3120
rect 3597 3116 3601 3120
rect 3619 3116 3623 3120
rect 3665 3116 3669 3120
rect 3673 3116 3677 3120
rect 3693 3116 3697 3120
rect 3703 3116 3707 3120
rect 3725 3116 3729 3120
rect 3771 3116 3775 3120
rect 3791 3116 3795 3120
rect 3865 3116 3869 3120
rect 3885 3116 3889 3120
rect 3905 3116 3909 3120
rect 3965 3116 3969 3120
rect 3985 3116 3989 3120
rect 4005 3116 4009 3120
rect 4051 3116 4055 3120
rect 4071 3116 4075 3120
rect 4091 3116 4095 3120
rect 4151 3116 4155 3120
rect 4171 3116 4175 3120
rect 4191 3116 4195 3120
rect 4251 3116 4255 3120
rect 4312 3116 4316 3120
rect 4320 3116 4324 3120
rect 4328 3116 4332 3120
rect 4411 3116 4415 3120
rect 4433 3116 4437 3120
rect 4443 3116 4447 3120
rect 4463 3116 4467 3120
rect 4471 3116 4475 3120
rect 4517 3116 4521 3120
rect 4539 3116 4543 3120
rect 4549 3116 4553 3120
rect 4571 3116 4575 3120
rect 4581 3116 4585 3120
rect 4601 3116 4605 3120
rect 4651 3116 4655 3120
rect 4671 3116 4675 3120
rect 4691 3116 4695 3120
rect 66 3071 70 3076
rect 40 3067 70 3071
rect 40 3019 46 3067
rect 74 3062 78 3076
rect 65 3055 78 3062
rect 65 3053 69 3055
rect 94 3053 98 3076
rect 102 3068 106 3076
rect 175 3070 179 3076
rect 102 3061 119 3068
rect 67 3041 69 3053
rect 46 3007 49 3019
rect 45 2984 49 3007
rect 65 2984 69 3041
rect 94 3012 98 3041
rect 113 3019 119 3061
rect 161 3058 173 3070
rect 85 3006 98 3012
rect 105 3007 113 3012
rect 105 3006 125 3007
rect 85 2984 89 3006
rect 105 2984 109 3006
rect 161 2984 165 3058
rect 195 3033 199 3076
rect 186 3021 199 3033
rect 183 2944 187 3021
rect 205 3019 209 3076
rect 205 3007 214 3019
rect 251 3008 255 3076
rect 273 3047 277 3096
rect 283 3075 287 3096
rect 303 3084 307 3096
rect 311 3092 315 3096
rect 311 3088 345 3092
rect 303 3080 333 3084
rect 303 3079 321 3080
rect 283 3071 307 3075
rect 205 2944 209 3007
rect 251 2996 253 3008
rect 251 2984 255 2996
rect 273 2989 277 3035
rect 269 2983 277 2989
rect 269 2954 273 2983
rect 301 2976 307 3071
rect 269 2947 277 2954
rect 273 2924 277 2947
rect 281 2924 285 2964
rect 301 2944 305 2976
rect 341 2962 345 3088
rect 357 2982 361 3096
rect 379 3084 383 3096
rect 381 3072 383 3084
rect 389 3084 393 3096
rect 389 3072 391 3084
rect 309 2950 333 2952
rect 309 2948 345 2950
rect 309 2944 313 2948
rect 355 2944 359 2970
rect 373 2962 377 3072
rect 411 3064 415 3096
rect 382 3060 415 3064
rect 382 2996 386 3060
rect 402 3011 406 3040
rect 421 3038 425 3096
rect 441 3039 445 3076
rect 491 3071 495 3076
rect 482 3064 495 3071
rect 402 3003 411 3011
rect 382 2984 385 2996
rect 375 2944 379 2950
rect 387 2944 391 2984
rect 407 2944 411 3003
rect 421 2944 425 3026
rect 441 2984 445 3027
rect 482 3019 486 3064
rect 511 3053 515 3076
rect 506 3041 515 3053
rect 482 2996 486 3007
rect 482 2988 500 2996
rect 496 2984 500 2988
rect 504 2984 508 3041
rect 531 2999 535 3076
rect 593 3056 597 3076
rect 589 3049 597 3056
rect 603 3056 607 3076
rect 693 3056 697 3076
rect 603 3049 617 3056
rect 589 3033 595 3049
rect 586 3021 595 3033
rect 526 2987 533 2999
rect 526 2944 530 2987
rect 591 2944 595 3021
rect 611 3033 617 3049
rect 683 3049 697 3056
rect 703 3056 707 3076
rect 703 3049 711 3056
rect 683 3033 689 3049
rect 611 3021 614 3033
rect 686 3021 689 3033
rect 611 2944 615 3021
rect 685 2944 689 3021
rect 705 3033 711 3049
rect 705 3021 714 3033
rect 705 2944 709 3021
rect 765 3019 769 3096
rect 785 3019 789 3096
rect 833 3056 837 3076
rect 829 3049 837 3056
rect 843 3056 847 3076
rect 843 3049 857 3056
rect 829 3033 835 3049
rect 826 3021 835 3033
rect 766 3007 781 3019
rect 777 2984 781 3007
rect 785 3007 794 3019
rect 785 2984 789 3007
rect 831 2944 835 3021
rect 851 3033 857 3049
rect 851 3021 854 3033
rect 851 2944 855 3021
rect 925 2999 929 3076
rect 945 3053 949 3076
rect 965 3071 969 3076
rect 965 3064 978 3071
rect 945 3041 954 3053
rect 927 2987 934 2999
rect 930 2944 934 2987
rect 952 2984 956 3041
rect 974 3019 978 3064
rect 974 2996 978 3007
rect 1025 2999 1029 3076
rect 1045 3053 1049 3076
rect 1065 3071 1069 3076
rect 1065 3064 1078 3071
rect 1045 3041 1054 3053
rect 960 2988 978 2996
rect 960 2984 964 2988
rect 1027 2987 1034 2999
rect 1030 2944 1034 2987
rect 1052 2984 1056 3041
rect 1074 3019 1078 3064
rect 1125 3019 1129 3096
rect 1145 3019 1149 3096
rect 1126 3007 1141 3019
rect 1074 2996 1078 3007
rect 1060 2988 1078 2996
rect 1060 2984 1064 2988
rect 1137 2984 1141 3007
rect 1145 3007 1154 3019
rect 1145 2984 1149 3007
rect 1205 2999 1209 3076
rect 1225 3053 1229 3076
rect 1245 3071 1249 3076
rect 1245 3064 1258 3071
rect 1225 3041 1234 3053
rect 1207 2987 1214 2999
rect 1210 2944 1214 2987
rect 1232 2984 1236 3041
rect 1254 3019 1258 3064
rect 1293 3056 1297 3076
rect 1289 3049 1297 3056
rect 1303 3056 1307 3076
rect 1303 3049 1317 3056
rect 1289 3033 1295 3049
rect 1286 3021 1295 3033
rect 1254 2996 1258 3007
rect 1240 2988 1258 2996
rect 1240 2984 1244 2988
rect 1291 2944 1295 3021
rect 1311 3033 1317 3049
rect 1385 3053 1389 3076
rect 1433 3056 1437 3076
rect 1385 3041 1394 3053
rect 1429 3049 1437 3056
rect 1443 3056 1447 3076
rect 1513 3056 1517 3076
rect 1443 3049 1457 3056
rect 1311 3021 1314 3033
rect 1311 2944 1315 3021
rect 1385 2984 1389 3041
rect 1429 3033 1435 3049
rect 1426 3021 1435 3033
rect 1431 2944 1435 3021
rect 1451 3033 1457 3049
rect 1509 3049 1517 3056
rect 1523 3056 1527 3076
rect 1523 3049 1537 3056
rect 1509 3033 1515 3049
rect 1451 3021 1454 3033
rect 1506 3021 1515 3033
rect 1451 2944 1455 3021
rect 1511 2944 1515 3021
rect 1531 3033 1537 3049
rect 1531 3021 1534 3033
rect 1531 2944 1535 3021
rect 1591 3019 1595 3096
rect 1613 3070 1617 3076
rect 1671 3071 1675 3076
rect 1615 3058 1617 3070
rect 1662 3064 1675 3071
rect 1662 3019 1666 3064
rect 1691 3053 1695 3076
rect 1686 3041 1695 3053
rect 1586 3007 1595 3019
rect 1591 2944 1595 3007
rect 1615 2990 1617 3002
rect 1613 2984 1617 2990
rect 1662 2996 1666 3007
rect 1662 2988 1680 2996
rect 1676 2984 1680 2988
rect 1684 2984 1688 3041
rect 1711 2999 1715 3076
rect 1771 3071 1775 3076
rect 1762 3064 1775 3071
rect 1762 3019 1766 3064
rect 1791 3053 1795 3076
rect 1786 3041 1795 3053
rect 1706 2987 1713 2999
rect 1762 2996 1766 3007
rect 1762 2988 1780 2996
rect 1706 2944 1710 2987
rect 1776 2984 1780 2988
rect 1784 2984 1788 3041
rect 1811 2999 1815 3076
rect 1871 3019 1875 3096
rect 1891 3019 1895 3096
rect 1954 3072 1958 3076
rect 1939 3066 1958 3072
rect 1939 3053 1946 3066
rect 1866 3007 1875 3019
rect 1806 2987 1813 2999
rect 1806 2944 1810 2987
rect 1871 2984 1875 3007
rect 1879 3007 1894 3019
rect 1879 2984 1883 3007
rect 1939 3004 1946 3041
rect 1962 3039 1966 3076
rect 1984 3053 1988 3096
rect 1986 3041 1995 3053
rect 1960 3004 1966 3027
rect 1939 2998 1955 3004
rect 1960 2998 1975 3004
rect 1951 2984 1955 2998
rect 1971 2984 1975 2998
rect 1991 2984 1995 3041
rect 2051 3039 2055 3096
rect 2111 3071 2115 3076
rect 2046 3027 2055 3039
rect 2051 2944 2055 3027
rect 2102 3064 2115 3071
rect 2102 3019 2106 3064
rect 2131 3053 2135 3076
rect 2126 3041 2135 3053
rect 2102 2996 2106 3007
rect 2102 2988 2120 2996
rect 2116 2984 2120 2988
rect 2124 2984 2128 3041
rect 2151 2999 2155 3076
rect 2211 3019 2215 3096
rect 2231 3019 2235 3096
rect 2313 3056 2317 3076
rect 2303 3049 2317 3056
rect 2323 3056 2327 3076
rect 2371 3071 2375 3076
rect 2362 3064 2375 3071
rect 2323 3049 2331 3056
rect 2303 3033 2309 3049
rect 2306 3021 2309 3033
rect 2206 3007 2215 3019
rect 2146 2987 2153 2999
rect 2146 2944 2150 2987
rect 2211 2984 2215 3007
rect 2219 3007 2234 3019
rect 2219 2984 2223 3007
rect 2305 2944 2309 3021
rect 2325 3033 2331 3049
rect 2325 3021 2334 3033
rect 2325 2944 2329 3021
rect 2362 3019 2366 3064
rect 2391 3053 2395 3076
rect 2386 3041 2395 3053
rect 2362 2996 2366 3007
rect 2362 2988 2380 2996
rect 2376 2984 2380 2988
rect 2384 2984 2388 3041
rect 2411 2999 2415 3076
rect 2471 3039 2475 3096
rect 2531 3071 2535 3076
rect 2466 3027 2475 3039
rect 2406 2987 2413 2999
rect 2406 2944 2410 2987
rect 2471 2944 2475 3027
rect 2522 3064 2535 3071
rect 2522 3019 2526 3064
rect 2551 3053 2555 3076
rect 2546 3041 2555 3053
rect 2522 2996 2526 3007
rect 2522 2988 2540 2996
rect 2536 2984 2540 2988
rect 2544 2984 2548 3041
rect 2571 2999 2575 3076
rect 2631 3019 2635 3096
rect 2653 3070 2657 3076
rect 2655 3058 2657 3070
rect 2713 3056 2717 3076
rect 2709 3049 2717 3056
rect 2723 3056 2727 3076
rect 2723 3049 2737 3056
rect 2709 3033 2715 3049
rect 2706 3021 2715 3033
rect 2626 3007 2635 3019
rect 2566 2987 2573 2999
rect 2566 2944 2570 2987
rect 2631 2944 2635 3007
rect 2655 2990 2657 3002
rect 2653 2984 2657 2990
rect 2711 2944 2715 3021
rect 2731 3033 2737 3049
rect 2795 3039 2799 3076
rect 2731 3021 2734 3033
rect 2815 3038 2819 3096
rect 2825 3064 2829 3096
rect 2847 3084 2851 3096
rect 2849 3072 2851 3084
rect 2857 3084 2861 3096
rect 2857 3072 2859 3084
rect 2825 3060 2858 3064
rect 2731 2944 2735 3021
rect 2795 2984 2799 3027
rect 2815 2944 2819 3026
rect 2834 3011 2838 3040
rect 2829 3003 2838 3011
rect 2829 2944 2833 3003
rect 2854 2996 2858 3060
rect 2855 2984 2858 2996
rect 2849 2944 2853 2984
rect 2863 2962 2867 3072
rect 2879 2982 2883 3096
rect 2925 3092 2929 3096
rect 2895 3088 2929 3092
rect 2861 2944 2865 2950
rect 2881 2944 2885 2970
rect 2895 2962 2899 3088
rect 2933 3084 2937 3096
rect 2907 3080 2937 3084
rect 2919 3079 2937 3080
rect 2953 3075 2957 3096
rect 2933 3071 2957 3075
rect 2933 2976 2939 3071
rect 2963 3047 2967 3096
rect 2963 2989 2967 3035
rect 2985 3008 2989 3076
rect 3045 3019 3049 3096
rect 3065 3019 3069 3096
rect 3132 3053 3136 3096
rect 3125 3041 3134 3053
rect 2987 2996 2989 3008
rect 3046 3007 3061 3019
rect 2963 2983 2971 2989
rect 2985 2984 2989 2996
rect 3057 2984 3061 3007
rect 3065 3007 3074 3019
rect 3065 2984 3069 3007
rect 3125 2984 3129 3041
rect 3154 3039 3158 3076
rect 3162 3072 3166 3076
rect 3162 3066 3181 3072
rect 3174 3053 3181 3066
rect 3154 3004 3160 3027
rect 3174 3004 3181 3041
rect 3211 3019 3215 3096
rect 3231 3019 3235 3096
rect 3295 3039 3299 3076
rect 3315 3038 3319 3096
rect 3325 3064 3329 3096
rect 3347 3084 3351 3096
rect 3349 3072 3351 3084
rect 3357 3084 3361 3096
rect 3357 3072 3359 3084
rect 3325 3060 3358 3064
rect 3206 3007 3215 3019
rect 3145 2998 3160 3004
rect 3165 2998 3181 3004
rect 3145 2984 3149 2998
rect 3165 2984 3169 2998
rect 3211 2984 3215 3007
rect 3219 3007 3234 3019
rect 3219 2984 3223 3007
rect 3295 2984 3299 3027
rect 2907 2950 2931 2952
rect 2895 2948 2931 2950
rect 2927 2944 2931 2948
rect 2935 2944 2939 2976
rect 2955 2924 2959 2964
rect 2967 2954 2971 2983
rect 2963 2947 2971 2954
rect 2963 2924 2967 2947
rect 3315 2944 3319 3026
rect 3334 3011 3338 3040
rect 3329 3003 3338 3011
rect 3329 2944 3333 3003
rect 3354 2996 3358 3060
rect 3355 2984 3358 2996
rect 3349 2944 3353 2984
rect 3363 2962 3367 3072
rect 3379 2982 3383 3096
rect 3425 3092 3429 3096
rect 3395 3088 3429 3092
rect 3361 2944 3365 2950
rect 3381 2944 3385 2970
rect 3395 2962 3399 3088
rect 3433 3084 3437 3096
rect 3407 3080 3437 3084
rect 3419 3079 3437 3080
rect 3453 3075 3457 3096
rect 3433 3071 3457 3075
rect 3433 2976 3439 3071
rect 3463 3047 3467 3096
rect 3463 2989 3467 3035
rect 3485 3008 3489 3076
rect 3535 3039 3539 3076
rect 3555 3038 3559 3096
rect 3565 3064 3569 3096
rect 3587 3084 3591 3096
rect 3589 3072 3591 3084
rect 3597 3084 3601 3096
rect 3597 3072 3599 3084
rect 3565 3060 3598 3064
rect 3487 2996 3489 3008
rect 3463 2983 3471 2989
rect 3485 2984 3489 2996
rect 3535 2984 3539 3027
rect 3407 2950 3431 2952
rect 3395 2948 3431 2950
rect 3427 2944 3431 2948
rect 3435 2944 3439 2976
rect 3455 2924 3459 2964
rect 3467 2954 3471 2983
rect 3463 2947 3471 2954
rect 3463 2924 3467 2947
rect 3555 2944 3559 3026
rect 3574 3011 3578 3040
rect 3569 3003 3578 3011
rect 3569 2944 3573 3003
rect 3594 2996 3598 3060
rect 3595 2984 3598 2996
rect 3589 2944 3593 2984
rect 3603 2962 3607 3072
rect 3619 2982 3623 3096
rect 3665 3092 3669 3096
rect 3635 3088 3669 3092
rect 3601 2944 3605 2950
rect 3621 2944 3625 2970
rect 3635 2962 3639 3088
rect 3673 3084 3677 3096
rect 3647 3080 3677 3084
rect 3659 3079 3677 3080
rect 3693 3075 3697 3096
rect 3673 3071 3697 3075
rect 3673 2976 3679 3071
rect 3703 3047 3707 3096
rect 3703 2989 3707 3035
rect 3725 3008 3729 3076
rect 3771 3019 3775 3096
rect 3791 3019 3795 3096
rect 3727 2996 3729 3008
rect 3766 3007 3775 3019
rect 3703 2983 3711 2989
rect 3725 2984 3729 2996
rect 3771 2984 3775 3007
rect 3779 3007 3794 3019
rect 3779 2984 3783 3007
rect 3865 2999 3869 3076
rect 3885 3053 3889 3076
rect 3905 3071 3909 3076
rect 3905 3064 3918 3071
rect 3885 3041 3894 3053
rect 3867 2987 3874 2999
rect 3647 2950 3671 2952
rect 3635 2948 3671 2950
rect 3667 2944 3671 2948
rect 3675 2944 3679 2976
rect 3695 2924 3699 2964
rect 3707 2954 3711 2983
rect 3703 2947 3711 2954
rect 3703 2924 3707 2947
rect 3870 2944 3874 2987
rect 3892 2984 3896 3041
rect 3914 3019 3918 3064
rect 3914 2996 3918 3007
rect 3965 2999 3969 3076
rect 3985 3053 3989 3076
rect 4005 3071 4009 3076
rect 4051 3071 4055 3076
rect 4005 3064 4018 3071
rect 3985 3041 3994 3053
rect 3900 2988 3918 2996
rect 3900 2984 3904 2988
rect 3967 2987 3974 2999
rect 3970 2944 3974 2987
rect 3992 2984 3996 3041
rect 4014 3019 4018 3064
rect 4042 3064 4055 3071
rect 4042 3019 4046 3064
rect 4071 3053 4075 3076
rect 4066 3041 4075 3053
rect 4014 2996 4018 3007
rect 4000 2988 4018 2996
rect 4042 2996 4046 3007
rect 4042 2988 4060 2996
rect 4000 2984 4004 2988
rect 4056 2984 4060 2988
rect 4064 2984 4068 3041
rect 4091 2999 4095 3076
rect 4151 3071 4155 3076
rect 4142 3064 4155 3071
rect 4142 3019 4146 3064
rect 4171 3053 4175 3076
rect 4166 3041 4175 3053
rect 4086 2987 4093 2999
rect 4142 2996 4146 3007
rect 4142 2988 4160 2996
rect 4086 2944 4090 2987
rect 4156 2984 4160 2988
rect 4164 2984 4168 3041
rect 4191 2999 4195 3076
rect 4251 3039 4255 3096
rect 4246 3027 4255 3039
rect 4186 2987 4193 2999
rect 4186 2944 4190 2987
rect 4251 2944 4255 3027
rect 4312 2999 4316 3056
rect 4306 2987 4316 2999
rect 4300 2956 4306 2987
rect 4320 2979 4324 3056
rect 4328 2999 4332 3056
rect 4411 3008 4415 3076
rect 4433 3047 4437 3096
rect 4443 3075 4447 3096
rect 4463 3084 4467 3096
rect 4471 3092 4475 3096
rect 4471 3088 4505 3092
rect 4463 3080 4493 3084
rect 4463 3079 4481 3080
rect 4443 3071 4467 3075
rect 4328 2987 4335 2999
rect 4347 2987 4355 2999
rect 4320 2960 4326 2967
rect 4320 2956 4335 2960
rect 4300 2952 4315 2956
rect 4311 2944 4315 2952
rect 4331 2944 4335 2956
rect 4351 2944 4355 2987
rect 4411 2996 4413 3008
rect 4411 2984 4415 2996
rect 4433 2989 4437 3035
rect 4429 2983 4437 2989
rect 4429 2954 4433 2983
rect 4461 2976 4467 3071
rect 4429 2947 4437 2954
rect 4433 2924 4437 2947
rect 4441 2924 4445 2964
rect 4461 2944 4465 2976
rect 4501 2962 4505 3088
rect 4517 2982 4521 3096
rect 4539 3084 4543 3096
rect 4541 3072 4543 3084
rect 4549 3084 4553 3096
rect 4549 3072 4551 3084
rect 4469 2950 4493 2952
rect 4469 2948 4505 2950
rect 4469 2944 4473 2948
rect 4515 2944 4519 2970
rect 4533 2962 4537 3072
rect 4571 3064 4575 3096
rect 4542 3060 4575 3064
rect 4542 2996 4546 3060
rect 4562 3011 4566 3040
rect 4581 3038 4585 3096
rect 4601 3039 4605 3076
rect 4651 3071 4655 3076
rect 4642 3064 4655 3071
rect 4562 3003 4571 3011
rect 4542 2984 4545 2996
rect 4535 2944 4539 2950
rect 4547 2944 4551 2984
rect 4567 2944 4571 3003
rect 4581 2944 4585 3026
rect 4601 2984 4605 3027
rect 4642 3019 4646 3064
rect 4671 3053 4675 3076
rect 4666 3041 4675 3053
rect 4642 2996 4646 3007
rect 4642 2988 4660 2996
rect 4656 2984 4660 2988
rect 4664 2984 4668 3041
rect 4691 2999 4695 3076
rect 4686 2987 4693 2999
rect 4686 2944 4690 2987
rect 45 2900 49 2904
rect 65 2900 69 2904
rect 85 2900 89 2904
rect 105 2900 109 2904
rect 161 2900 165 2904
rect 183 2900 187 2904
rect 205 2900 209 2904
rect 251 2900 255 2904
rect 273 2900 277 2904
rect 281 2900 285 2904
rect 301 2900 305 2904
rect 309 2900 313 2904
rect 355 2900 359 2904
rect 375 2900 379 2904
rect 387 2900 391 2904
rect 407 2900 411 2904
rect 421 2900 425 2904
rect 441 2900 445 2904
rect 496 2900 500 2904
rect 504 2900 508 2904
rect 526 2900 530 2904
rect 591 2900 595 2904
rect 611 2900 615 2904
rect 685 2900 689 2904
rect 705 2900 709 2904
rect 777 2900 781 2904
rect 785 2900 789 2904
rect 831 2900 835 2904
rect 851 2900 855 2904
rect 930 2900 934 2904
rect 952 2900 956 2904
rect 960 2900 964 2904
rect 1030 2900 1034 2904
rect 1052 2900 1056 2904
rect 1060 2900 1064 2904
rect 1137 2900 1141 2904
rect 1145 2900 1149 2904
rect 1210 2900 1214 2904
rect 1232 2900 1236 2904
rect 1240 2900 1244 2904
rect 1291 2900 1295 2904
rect 1311 2900 1315 2904
rect 1385 2900 1389 2904
rect 1431 2900 1435 2904
rect 1451 2900 1455 2904
rect 1511 2900 1515 2904
rect 1531 2900 1535 2904
rect 1591 2900 1595 2904
rect 1613 2900 1617 2904
rect 1676 2900 1680 2904
rect 1684 2900 1688 2904
rect 1706 2900 1710 2904
rect 1776 2900 1780 2904
rect 1784 2900 1788 2904
rect 1806 2900 1810 2904
rect 1871 2900 1875 2904
rect 1879 2900 1883 2904
rect 1951 2900 1955 2904
rect 1971 2900 1975 2904
rect 1991 2900 1995 2904
rect 2051 2900 2055 2904
rect 2116 2900 2120 2904
rect 2124 2900 2128 2904
rect 2146 2900 2150 2904
rect 2211 2900 2215 2904
rect 2219 2900 2223 2904
rect 2305 2900 2309 2904
rect 2325 2900 2329 2904
rect 2376 2900 2380 2904
rect 2384 2900 2388 2904
rect 2406 2900 2410 2904
rect 2471 2900 2475 2904
rect 2536 2900 2540 2904
rect 2544 2900 2548 2904
rect 2566 2900 2570 2904
rect 2631 2900 2635 2904
rect 2653 2900 2657 2904
rect 2711 2900 2715 2904
rect 2731 2900 2735 2904
rect 2795 2900 2799 2904
rect 2815 2900 2819 2904
rect 2829 2900 2833 2904
rect 2849 2900 2853 2904
rect 2861 2900 2865 2904
rect 2881 2900 2885 2904
rect 2927 2900 2931 2904
rect 2935 2900 2939 2904
rect 2955 2900 2959 2904
rect 2963 2900 2967 2904
rect 2985 2900 2989 2904
rect 3057 2900 3061 2904
rect 3065 2900 3069 2904
rect 3125 2900 3129 2904
rect 3145 2900 3149 2904
rect 3165 2900 3169 2904
rect 3211 2900 3215 2904
rect 3219 2900 3223 2904
rect 3295 2900 3299 2904
rect 3315 2900 3319 2904
rect 3329 2900 3333 2904
rect 3349 2900 3353 2904
rect 3361 2900 3365 2904
rect 3381 2900 3385 2904
rect 3427 2900 3431 2904
rect 3435 2900 3439 2904
rect 3455 2900 3459 2904
rect 3463 2900 3467 2904
rect 3485 2900 3489 2904
rect 3535 2900 3539 2904
rect 3555 2900 3559 2904
rect 3569 2900 3573 2904
rect 3589 2900 3593 2904
rect 3601 2900 3605 2904
rect 3621 2900 3625 2904
rect 3667 2900 3671 2904
rect 3675 2900 3679 2904
rect 3695 2900 3699 2904
rect 3703 2900 3707 2904
rect 3725 2900 3729 2904
rect 3771 2900 3775 2904
rect 3779 2900 3783 2904
rect 3870 2900 3874 2904
rect 3892 2900 3896 2904
rect 3900 2900 3904 2904
rect 3970 2900 3974 2904
rect 3992 2900 3996 2904
rect 4000 2900 4004 2904
rect 4056 2900 4060 2904
rect 4064 2900 4068 2904
rect 4086 2900 4090 2904
rect 4156 2900 4160 2904
rect 4164 2900 4168 2904
rect 4186 2900 4190 2904
rect 4251 2900 4255 2904
rect 4311 2900 4315 2904
rect 4331 2900 4335 2904
rect 4351 2900 4355 2904
rect 4411 2900 4415 2904
rect 4433 2900 4437 2904
rect 4441 2900 4445 2904
rect 4461 2900 4465 2904
rect 4469 2900 4473 2904
rect 4515 2900 4519 2904
rect 4535 2900 4539 2904
rect 4547 2900 4551 2904
rect 4567 2900 4571 2904
rect 4581 2900 4585 2904
rect 4601 2900 4605 2904
rect 4656 2900 4660 2904
rect 4664 2900 4668 2904
rect 4686 2900 4690 2904
rect 45 2876 49 2880
rect 110 2876 114 2880
rect 132 2876 136 2880
rect 140 2876 144 2880
rect 191 2876 195 2880
rect 211 2876 215 2880
rect 231 2876 235 2880
rect 251 2876 255 2880
rect 311 2876 315 2880
rect 331 2876 335 2880
rect 391 2876 395 2880
rect 413 2876 417 2880
rect 435 2876 439 2880
rect 510 2876 514 2880
rect 532 2876 536 2880
rect 540 2876 544 2880
rect 591 2876 595 2880
rect 611 2876 615 2880
rect 685 2876 689 2880
rect 745 2876 749 2880
rect 791 2876 795 2880
rect 811 2876 815 2880
rect 871 2876 875 2880
rect 893 2876 897 2880
rect 915 2876 919 2880
rect 990 2876 994 2880
rect 1012 2876 1016 2880
rect 1020 2876 1024 2880
rect 1071 2876 1075 2880
rect 1091 2876 1095 2880
rect 1170 2876 1174 2880
rect 1192 2876 1196 2880
rect 1200 2876 1204 2880
rect 1251 2876 1255 2880
rect 1273 2876 1277 2880
rect 1281 2876 1285 2880
rect 1301 2876 1305 2880
rect 1309 2876 1313 2880
rect 1355 2876 1359 2880
rect 1375 2876 1379 2880
rect 1387 2876 1391 2880
rect 1407 2876 1411 2880
rect 1421 2876 1425 2880
rect 1441 2876 1445 2880
rect 1503 2876 1507 2880
rect 1525 2876 1529 2880
rect 1575 2876 1579 2880
rect 1595 2876 1599 2880
rect 1609 2876 1613 2880
rect 1629 2876 1633 2880
rect 1641 2876 1645 2880
rect 1661 2876 1665 2880
rect 1707 2876 1711 2880
rect 1715 2876 1719 2880
rect 1735 2876 1739 2880
rect 1743 2876 1747 2880
rect 1765 2876 1769 2880
rect 1816 2876 1820 2880
rect 1824 2876 1828 2880
rect 1846 2876 1850 2880
rect 1911 2876 1915 2880
rect 1971 2876 1975 2880
rect 1981 2876 1985 2880
rect 2011 2876 2015 2880
rect 2021 2876 2025 2880
rect 2117 2876 2121 2880
rect 2125 2876 2129 2880
rect 2197 2876 2201 2880
rect 2205 2876 2209 2880
rect 2277 2876 2281 2880
rect 2285 2876 2289 2880
rect 2331 2876 2335 2880
rect 2417 2876 2421 2880
rect 2425 2876 2429 2880
rect 2471 2876 2475 2880
rect 2531 2876 2535 2880
rect 2553 2876 2557 2880
rect 2575 2876 2579 2880
rect 2636 2876 2640 2880
rect 2644 2876 2648 2880
rect 2666 2876 2670 2880
rect 2736 2876 2740 2880
rect 2744 2876 2748 2880
rect 2766 2876 2770 2880
rect 2831 2876 2835 2880
rect 2851 2876 2855 2880
rect 2915 2876 2919 2880
rect 2935 2876 2939 2880
rect 2949 2876 2953 2880
rect 2969 2876 2973 2880
rect 2981 2876 2985 2880
rect 3001 2876 3005 2880
rect 3047 2876 3051 2880
rect 3055 2876 3059 2880
rect 3075 2876 3079 2880
rect 3083 2876 3087 2880
rect 3105 2876 3109 2880
rect 3155 2876 3159 2880
rect 3175 2876 3179 2880
rect 3189 2876 3193 2880
rect 3209 2876 3213 2880
rect 3221 2876 3225 2880
rect 3241 2876 3245 2880
rect 3287 2876 3291 2880
rect 3295 2876 3299 2880
rect 3315 2876 3319 2880
rect 3323 2876 3327 2880
rect 3345 2876 3349 2880
rect 3405 2876 3409 2880
rect 3477 2876 3481 2880
rect 3485 2876 3489 2880
rect 3545 2876 3549 2880
rect 3595 2876 3599 2880
rect 3615 2876 3619 2880
rect 3629 2876 3633 2880
rect 3649 2876 3653 2880
rect 3661 2876 3665 2880
rect 3681 2876 3685 2880
rect 3727 2876 3731 2880
rect 3735 2876 3739 2880
rect 3755 2876 3759 2880
rect 3763 2876 3767 2880
rect 3785 2876 3789 2880
rect 3845 2876 3849 2880
rect 3865 2876 3869 2880
rect 3885 2876 3889 2880
rect 3905 2876 3909 2880
rect 3977 2876 3981 2880
rect 3985 2876 3989 2880
rect 4036 2876 4040 2880
rect 4044 2876 4048 2880
rect 4066 2876 4070 2880
rect 4150 2876 4154 2880
rect 4172 2876 4176 2880
rect 4180 2876 4184 2880
rect 4231 2876 4235 2880
rect 4239 2876 4243 2880
rect 4315 2876 4319 2880
rect 4335 2876 4339 2880
rect 4349 2876 4353 2880
rect 4369 2876 4373 2880
rect 4381 2876 4385 2880
rect 4401 2876 4405 2880
rect 4447 2876 4451 2880
rect 4455 2876 4459 2880
rect 4475 2876 4479 2880
rect 4483 2876 4487 2880
rect 4505 2876 4509 2880
rect 4556 2876 4560 2880
rect 4564 2876 4568 2880
rect 4586 2876 4590 2880
rect 4651 2876 4655 2880
rect 4671 2876 4675 2880
rect 45 2753 49 2836
rect 110 2793 114 2836
rect 107 2781 114 2793
rect 45 2741 54 2753
rect 45 2684 49 2741
rect 105 2704 109 2781
rect 132 2739 136 2796
rect 140 2792 144 2796
rect 140 2784 158 2792
rect 154 2773 158 2784
rect 191 2774 195 2796
rect 211 2774 215 2796
rect 175 2773 195 2774
rect 187 2768 195 2773
rect 202 2768 215 2774
rect 125 2727 134 2739
rect 125 2704 129 2727
rect 154 2716 158 2761
rect 145 2709 158 2716
rect 181 2719 187 2761
rect 202 2739 206 2768
rect 231 2739 235 2796
rect 251 2773 255 2796
rect 251 2761 254 2773
rect 231 2727 233 2739
rect 181 2712 198 2719
rect 145 2704 149 2709
rect 194 2704 198 2712
rect 202 2704 206 2727
rect 231 2725 235 2727
rect 222 2718 235 2725
rect 222 2704 226 2718
rect 254 2713 260 2761
rect 311 2759 315 2836
rect 306 2747 315 2759
rect 309 2731 315 2747
rect 331 2759 335 2836
rect 391 2773 395 2836
rect 386 2761 395 2773
rect 331 2747 334 2759
rect 331 2731 337 2747
rect 309 2724 317 2731
rect 230 2709 260 2713
rect 230 2704 234 2709
rect 313 2704 317 2724
rect 323 2724 337 2731
rect 323 2704 327 2724
rect 391 2704 395 2761
rect 413 2759 417 2836
rect 401 2747 414 2759
rect 401 2704 405 2747
rect 435 2722 439 2796
rect 510 2793 514 2836
rect 507 2781 514 2793
rect 427 2710 439 2722
rect 421 2704 425 2710
rect 505 2704 509 2781
rect 532 2739 536 2796
rect 540 2792 544 2796
rect 540 2784 558 2792
rect 554 2773 558 2784
rect 525 2727 534 2739
rect 525 2704 529 2727
rect 554 2716 558 2761
rect 591 2759 595 2836
rect 586 2747 595 2759
rect 589 2731 595 2747
rect 611 2759 615 2836
rect 611 2747 614 2759
rect 611 2731 617 2747
rect 589 2724 597 2731
rect 545 2709 558 2716
rect 545 2704 549 2709
rect 593 2704 597 2724
rect 603 2724 617 2731
rect 685 2739 689 2796
rect 745 2739 749 2796
rect 791 2759 795 2836
rect 786 2747 795 2759
rect 685 2727 694 2739
rect 745 2727 754 2739
rect 789 2731 795 2747
rect 811 2759 815 2836
rect 871 2773 875 2836
rect 866 2761 875 2773
rect 811 2747 814 2759
rect 811 2731 817 2747
rect 603 2704 607 2724
rect 685 2704 689 2727
rect 745 2704 749 2727
rect 789 2724 797 2731
rect 793 2704 797 2724
rect 803 2724 817 2731
rect 803 2704 807 2724
rect 871 2704 875 2761
rect 893 2759 897 2836
rect 881 2747 894 2759
rect 881 2704 885 2747
rect 915 2722 919 2796
rect 990 2793 994 2836
rect 987 2781 994 2793
rect 907 2710 919 2722
rect 901 2704 905 2710
rect 985 2704 989 2781
rect 1012 2739 1016 2796
rect 1020 2792 1024 2796
rect 1020 2784 1038 2792
rect 1034 2773 1038 2784
rect 1005 2727 1014 2739
rect 1005 2704 1009 2727
rect 1034 2716 1038 2761
rect 1071 2759 1075 2836
rect 1066 2747 1075 2759
rect 1069 2731 1075 2747
rect 1091 2759 1095 2836
rect 1170 2793 1174 2836
rect 1273 2833 1277 2856
rect 1269 2826 1277 2833
rect 1269 2797 1273 2826
rect 1281 2816 1285 2856
rect 1301 2804 1305 2836
rect 1309 2832 1313 2836
rect 1309 2830 1345 2832
rect 1309 2828 1333 2830
rect 1167 2781 1174 2793
rect 1091 2747 1094 2759
rect 1091 2731 1097 2747
rect 1069 2724 1077 2731
rect 1025 2709 1038 2716
rect 1025 2704 1029 2709
rect 1073 2704 1077 2724
rect 1083 2724 1097 2731
rect 1083 2704 1087 2724
rect 1165 2704 1169 2781
rect 1192 2739 1196 2796
rect 1200 2792 1204 2796
rect 1200 2784 1218 2792
rect 1214 2773 1218 2784
rect 1251 2784 1255 2796
rect 1269 2791 1277 2797
rect 1251 2772 1253 2784
rect 1185 2727 1194 2739
rect 1185 2704 1189 2727
rect 1214 2716 1218 2761
rect 1205 2709 1218 2716
rect 1205 2704 1209 2709
rect 1251 2704 1255 2772
rect 1273 2745 1277 2791
rect 1273 2684 1277 2733
rect 1301 2709 1307 2804
rect 1283 2705 1307 2709
rect 1283 2684 1287 2705
rect 1303 2700 1321 2701
rect 1303 2696 1333 2700
rect 1303 2684 1307 2696
rect 1341 2692 1345 2818
rect 1355 2810 1359 2836
rect 1375 2830 1379 2836
rect 1311 2688 1345 2692
rect 1311 2684 1315 2688
rect 1357 2684 1361 2798
rect 1373 2708 1377 2818
rect 1387 2796 1391 2836
rect 1382 2784 1385 2796
rect 1382 2720 1386 2784
rect 1407 2777 1411 2836
rect 1402 2769 1411 2777
rect 1402 2740 1406 2769
rect 1421 2754 1425 2836
rect 1441 2753 1445 2796
rect 1503 2790 1507 2796
rect 1503 2778 1505 2790
rect 1525 2773 1529 2836
rect 1525 2761 1534 2773
rect 1382 2716 1415 2720
rect 1381 2696 1383 2708
rect 1379 2684 1383 2696
rect 1389 2696 1391 2708
rect 1389 2684 1393 2696
rect 1411 2684 1415 2716
rect 1421 2684 1425 2742
rect 1441 2704 1445 2741
rect 1503 2710 1505 2722
rect 1503 2704 1507 2710
rect 1525 2684 1529 2761
rect 1575 2753 1579 2796
rect 1595 2754 1599 2836
rect 1609 2777 1613 2836
rect 1629 2796 1633 2836
rect 1641 2830 1645 2836
rect 1635 2784 1638 2796
rect 1609 2769 1618 2777
rect 1575 2704 1579 2741
rect 1595 2684 1599 2742
rect 1614 2740 1618 2769
rect 1634 2720 1638 2784
rect 1605 2716 1638 2720
rect 1605 2684 1609 2716
rect 1643 2708 1647 2818
rect 1661 2810 1665 2836
rect 1707 2832 1711 2836
rect 1675 2830 1711 2832
rect 1687 2828 1711 2830
rect 1629 2696 1631 2708
rect 1627 2684 1631 2696
rect 1637 2696 1639 2708
rect 1637 2684 1641 2696
rect 1659 2684 1663 2798
rect 1675 2692 1679 2818
rect 1715 2804 1719 2836
rect 1735 2816 1739 2856
rect 1743 2833 1747 2856
rect 1743 2826 1751 2833
rect 1713 2709 1719 2804
rect 1747 2797 1751 2826
rect 1743 2791 1751 2797
rect 1743 2745 1747 2791
rect 1765 2784 1769 2796
rect 1816 2792 1820 2796
rect 1767 2772 1769 2784
rect 1802 2784 1820 2792
rect 1802 2773 1806 2784
rect 1713 2705 1737 2709
rect 1699 2700 1717 2701
rect 1687 2696 1717 2700
rect 1675 2688 1709 2692
rect 1705 2684 1709 2688
rect 1713 2684 1717 2696
rect 1733 2684 1737 2705
rect 1743 2684 1747 2733
rect 1765 2704 1769 2772
rect 1802 2716 1806 2761
rect 1824 2739 1828 2796
rect 1846 2793 1850 2836
rect 1846 2781 1853 2793
rect 1826 2727 1835 2739
rect 1802 2709 1815 2716
rect 1811 2704 1815 2709
rect 1831 2704 1835 2727
rect 1851 2704 1855 2781
rect 1911 2753 1915 2836
rect 1971 2792 1975 2796
rect 1961 2788 1975 2792
rect 1981 2792 1985 2796
rect 1981 2788 1995 2792
rect 1961 2773 1966 2788
rect 1906 2741 1915 2753
rect 1911 2684 1915 2741
rect 1960 2715 1966 2761
rect 1989 2739 1995 2788
rect 2011 2739 2015 2796
rect 2021 2792 2025 2796
rect 2021 2788 2035 2792
rect 2031 2773 2035 2788
rect 2117 2773 2121 2796
rect 2031 2761 2033 2773
rect 2106 2761 2121 2773
rect 2125 2773 2129 2796
rect 2197 2773 2201 2796
rect 2125 2761 2134 2773
rect 2186 2761 2201 2773
rect 2205 2773 2209 2796
rect 2277 2773 2281 2796
rect 2205 2761 2214 2773
rect 2266 2761 2281 2773
rect 2285 2773 2289 2796
rect 2285 2761 2294 2773
rect 1986 2727 1995 2739
rect 1960 2711 1975 2715
rect 1971 2704 1975 2711
rect 1991 2704 1995 2727
rect 2011 2704 2015 2727
rect 2031 2704 2035 2761
rect 2105 2684 2109 2761
rect 2125 2684 2129 2761
rect 2185 2684 2189 2761
rect 2205 2684 2209 2761
rect 2265 2684 2269 2761
rect 2285 2684 2289 2761
rect 2331 2753 2335 2836
rect 2417 2773 2421 2796
rect 2406 2761 2421 2773
rect 2425 2773 2429 2796
rect 2425 2761 2434 2773
rect 2326 2741 2335 2753
rect 2331 2684 2335 2741
rect 2405 2684 2409 2761
rect 2425 2684 2429 2761
rect 2471 2753 2475 2836
rect 2531 2773 2535 2836
rect 2526 2761 2535 2773
rect 2466 2741 2475 2753
rect 2471 2684 2475 2741
rect 2531 2704 2535 2761
rect 2553 2759 2557 2836
rect 2541 2747 2554 2759
rect 2541 2704 2545 2747
rect 2575 2722 2579 2796
rect 2636 2792 2640 2796
rect 2622 2784 2640 2792
rect 2622 2773 2626 2784
rect 2567 2710 2579 2722
rect 2622 2716 2626 2761
rect 2644 2739 2648 2796
rect 2666 2793 2670 2836
rect 2666 2781 2673 2793
rect 2736 2792 2740 2796
rect 2722 2784 2740 2792
rect 2646 2727 2655 2739
rect 2561 2704 2565 2710
rect 2622 2709 2635 2716
rect 2631 2704 2635 2709
rect 2651 2704 2655 2727
rect 2671 2704 2675 2781
rect 2722 2773 2726 2784
rect 2722 2716 2726 2761
rect 2744 2739 2748 2796
rect 2766 2793 2770 2836
rect 2766 2781 2773 2793
rect 2746 2727 2755 2739
rect 2722 2709 2735 2716
rect 2731 2704 2735 2709
rect 2751 2704 2755 2727
rect 2771 2704 2775 2781
rect 2831 2759 2835 2836
rect 2826 2747 2835 2759
rect 2829 2731 2835 2747
rect 2851 2759 2855 2836
rect 2851 2747 2854 2759
rect 2915 2753 2919 2796
rect 2935 2754 2939 2836
rect 2949 2777 2953 2836
rect 2969 2796 2973 2836
rect 2981 2830 2985 2836
rect 2975 2784 2978 2796
rect 2949 2769 2958 2777
rect 2851 2731 2857 2747
rect 2829 2724 2837 2731
rect 2833 2704 2837 2724
rect 2843 2724 2857 2731
rect 2843 2704 2847 2724
rect 2915 2704 2919 2741
rect 2935 2684 2939 2742
rect 2954 2740 2958 2769
rect 2974 2720 2978 2784
rect 2945 2716 2978 2720
rect 2945 2684 2949 2716
rect 2983 2708 2987 2818
rect 3001 2810 3005 2836
rect 3047 2832 3051 2836
rect 3015 2830 3051 2832
rect 3027 2828 3051 2830
rect 2969 2696 2971 2708
rect 2967 2684 2971 2696
rect 2977 2696 2979 2708
rect 2977 2684 2981 2696
rect 2999 2684 3003 2798
rect 3015 2692 3019 2818
rect 3055 2804 3059 2836
rect 3075 2816 3079 2856
rect 3083 2833 3087 2856
rect 3083 2826 3091 2833
rect 3053 2709 3059 2804
rect 3087 2797 3091 2826
rect 3083 2791 3091 2797
rect 3083 2745 3087 2791
rect 3105 2784 3109 2796
rect 3107 2772 3109 2784
rect 3053 2705 3077 2709
rect 3039 2700 3057 2701
rect 3027 2696 3057 2700
rect 3015 2688 3049 2692
rect 3045 2684 3049 2688
rect 3053 2684 3057 2696
rect 3073 2684 3077 2705
rect 3083 2684 3087 2733
rect 3105 2704 3109 2772
rect 3155 2753 3159 2796
rect 3175 2754 3179 2836
rect 3189 2777 3193 2836
rect 3209 2796 3213 2836
rect 3221 2830 3225 2836
rect 3215 2784 3218 2796
rect 3189 2769 3198 2777
rect 3155 2704 3159 2741
rect 3175 2684 3179 2742
rect 3194 2740 3198 2769
rect 3214 2720 3218 2784
rect 3185 2716 3218 2720
rect 3185 2684 3189 2716
rect 3223 2708 3227 2818
rect 3241 2810 3245 2836
rect 3287 2832 3291 2836
rect 3255 2830 3291 2832
rect 3267 2828 3291 2830
rect 3209 2696 3211 2708
rect 3207 2684 3211 2696
rect 3217 2696 3219 2708
rect 3217 2684 3221 2696
rect 3239 2684 3243 2798
rect 3255 2692 3259 2818
rect 3295 2804 3299 2836
rect 3315 2816 3319 2856
rect 3323 2833 3327 2856
rect 3323 2826 3331 2833
rect 3293 2709 3299 2804
rect 3327 2797 3331 2826
rect 3323 2791 3331 2797
rect 3323 2745 3327 2791
rect 3345 2784 3349 2796
rect 3347 2772 3349 2784
rect 3293 2705 3317 2709
rect 3279 2700 3297 2701
rect 3267 2696 3297 2700
rect 3255 2688 3289 2692
rect 3285 2684 3289 2688
rect 3293 2684 3297 2696
rect 3313 2684 3317 2705
rect 3323 2684 3327 2733
rect 3345 2704 3349 2772
rect 3405 2753 3409 2836
rect 3477 2773 3481 2796
rect 3466 2761 3481 2773
rect 3485 2773 3489 2796
rect 3485 2761 3494 2773
rect 3405 2741 3414 2753
rect 3405 2684 3409 2741
rect 3465 2684 3469 2761
rect 3485 2684 3489 2761
rect 3545 2739 3549 2796
rect 3595 2753 3599 2796
rect 3615 2754 3619 2836
rect 3629 2777 3633 2836
rect 3649 2796 3653 2836
rect 3661 2830 3665 2836
rect 3655 2784 3658 2796
rect 3629 2769 3638 2777
rect 3545 2727 3554 2739
rect 3545 2704 3549 2727
rect 3595 2704 3599 2741
rect 3615 2684 3619 2742
rect 3634 2740 3638 2769
rect 3654 2720 3658 2784
rect 3625 2716 3658 2720
rect 3625 2684 3629 2716
rect 3663 2708 3667 2818
rect 3681 2810 3685 2836
rect 3727 2832 3731 2836
rect 3695 2830 3731 2832
rect 3707 2828 3731 2830
rect 3649 2696 3651 2708
rect 3647 2684 3651 2696
rect 3657 2696 3659 2708
rect 3657 2684 3661 2696
rect 3679 2684 3683 2798
rect 3695 2692 3699 2818
rect 3735 2804 3739 2836
rect 3755 2816 3759 2856
rect 3763 2833 3767 2856
rect 3763 2826 3771 2833
rect 3733 2709 3739 2804
rect 3767 2797 3771 2826
rect 3763 2791 3771 2797
rect 3763 2745 3767 2791
rect 3785 2784 3789 2796
rect 3787 2772 3789 2784
rect 3845 2773 3849 2796
rect 3733 2705 3757 2709
rect 3719 2700 3737 2701
rect 3707 2696 3737 2700
rect 3695 2688 3729 2692
rect 3725 2684 3729 2688
rect 3733 2684 3737 2696
rect 3753 2684 3757 2705
rect 3763 2684 3767 2733
rect 3785 2704 3789 2772
rect 3846 2761 3849 2773
rect 3840 2713 3846 2761
rect 3865 2739 3869 2796
rect 3885 2774 3889 2796
rect 3905 2774 3909 2796
rect 3885 2768 3898 2774
rect 3905 2773 3925 2774
rect 3977 2773 3981 2796
rect 3905 2768 3913 2773
rect 3894 2739 3898 2768
rect 3966 2761 3981 2773
rect 3985 2773 3989 2796
rect 4036 2792 4040 2796
rect 4022 2784 4040 2792
rect 4022 2773 4026 2784
rect 3985 2761 3994 2773
rect 3867 2727 3869 2739
rect 3865 2725 3869 2727
rect 3865 2718 3878 2725
rect 3840 2709 3870 2713
rect 3866 2704 3870 2709
rect 3874 2704 3878 2718
rect 3894 2704 3898 2727
rect 3913 2719 3919 2761
rect 3902 2712 3919 2719
rect 3902 2704 3906 2712
rect 3965 2684 3969 2761
rect 3985 2684 3989 2761
rect 4022 2716 4026 2761
rect 4044 2739 4048 2796
rect 4066 2793 4070 2836
rect 4150 2793 4154 2836
rect 4066 2781 4073 2793
rect 4147 2781 4154 2793
rect 4046 2727 4055 2739
rect 4022 2709 4035 2716
rect 4031 2704 4035 2709
rect 4051 2704 4055 2727
rect 4071 2704 4075 2781
rect 4145 2704 4149 2781
rect 4172 2739 4176 2796
rect 4180 2792 4184 2796
rect 4180 2784 4198 2792
rect 4194 2773 4198 2784
rect 4231 2773 4235 2796
rect 4226 2761 4235 2773
rect 4239 2773 4243 2796
rect 4239 2761 4254 2773
rect 4165 2727 4174 2739
rect 4165 2704 4169 2727
rect 4194 2716 4198 2761
rect 4185 2709 4198 2716
rect 4185 2704 4189 2709
rect 4231 2684 4235 2761
rect 4251 2684 4255 2761
rect 4315 2753 4319 2796
rect 4335 2754 4339 2836
rect 4349 2777 4353 2836
rect 4369 2796 4373 2836
rect 4381 2830 4385 2836
rect 4375 2784 4378 2796
rect 4349 2769 4358 2777
rect 4315 2704 4319 2741
rect 4335 2684 4339 2742
rect 4354 2740 4358 2769
rect 4374 2720 4378 2784
rect 4345 2716 4378 2720
rect 4345 2684 4349 2716
rect 4383 2708 4387 2818
rect 4401 2810 4405 2836
rect 4447 2832 4451 2836
rect 4415 2830 4451 2832
rect 4427 2828 4451 2830
rect 4369 2696 4371 2708
rect 4367 2684 4371 2696
rect 4377 2696 4379 2708
rect 4377 2684 4381 2696
rect 4399 2684 4403 2798
rect 4415 2692 4419 2818
rect 4455 2804 4459 2836
rect 4475 2816 4479 2856
rect 4483 2833 4487 2856
rect 4483 2826 4491 2833
rect 4453 2709 4459 2804
rect 4487 2797 4491 2826
rect 4483 2791 4491 2797
rect 4483 2745 4487 2791
rect 4505 2784 4509 2796
rect 4556 2792 4560 2796
rect 4507 2772 4509 2784
rect 4542 2784 4560 2792
rect 4542 2773 4546 2784
rect 4453 2705 4477 2709
rect 4439 2700 4457 2701
rect 4427 2696 4457 2700
rect 4415 2688 4449 2692
rect 4445 2684 4449 2688
rect 4453 2684 4457 2696
rect 4473 2684 4477 2705
rect 4483 2684 4487 2733
rect 4505 2704 4509 2772
rect 4542 2716 4546 2761
rect 4564 2739 4568 2796
rect 4586 2793 4590 2836
rect 4586 2781 4593 2793
rect 4566 2727 4575 2739
rect 4542 2709 4555 2716
rect 4551 2704 4555 2709
rect 4571 2704 4575 2727
rect 4591 2704 4595 2781
rect 4651 2759 4655 2836
rect 4646 2747 4655 2759
rect 4649 2731 4655 2747
rect 4671 2759 4675 2836
rect 4671 2747 4674 2759
rect 4671 2731 4677 2747
rect 4649 2724 4657 2731
rect 4653 2704 4657 2724
rect 4663 2724 4677 2731
rect 4663 2704 4667 2724
rect 45 2660 49 2664
rect 105 2660 109 2664
rect 125 2660 129 2664
rect 145 2660 149 2664
rect 194 2660 198 2664
rect 202 2660 206 2664
rect 222 2660 226 2664
rect 230 2660 234 2664
rect 313 2660 317 2664
rect 323 2660 327 2664
rect 391 2660 395 2664
rect 401 2660 405 2664
rect 421 2660 425 2664
rect 505 2660 509 2664
rect 525 2660 529 2664
rect 545 2660 549 2664
rect 593 2660 597 2664
rect 603 2660 607 2664
rect 685 2660 689 2664
rect 745 2660 749 2664
rect 793 2660 797 2664
rect 803 2660 807 2664
rect 871 2660 875 2664
rect 881 2660 885 2664
rect 901 2660 905 2664
rect 985 2660 989 2664
rect 1005 2660 1009 2664
rect 1025 2660 1029 2664
rect 1073 2660 1077 2664
rect 1083 2660 1087 2664
rect 1165 2660 1169 2664
rect 1185 2660 1189 2664
rect 1205 2660 1209 2664
rect 1251 2660 1255 2664
rect 1273 2660 1277 2664
rect 1283 2660 1287 2664
rect 1303 2660 1307 2664
rect 1311 2660 1315 2664
rect 1357 2660 1361 2664
rect 1379 2660 1383 2664
rect 1389 2660 1393 2664
rect 1411 2660 1415 2664
rect 1421 2660 1425 2664
rect 1441 2660 1445 2664
rect 1503 2660 1507 2664
rect 1525 2660 1529 2664
rect 1575 2660 1579 2664
rect 1595 2660 1599 2664
rect 1605 2660 1609 2664
rect 1627 2660 1631 2664
rect 1637 2660 1641 2664
rect 1659 2660 1663 2664
rect 1705 2660 1709 2664
rect 1713 2660 1717 2664
rect 1733 2660 1737 2664
rect 1743 2660 1747 2664
rect 1765 2660 1769 2664
rect 1811 2660 1815 2664
rect 1831 2660 1835 2664
rect 1851 2660 1855 2664
rect 1911 2660 1915 2664
rect 1971 2660 1975 2664
rect 1991 2660 1995 2664
rect 2011 2660 2015 2664
rect 2031 2660 2035 2664
rect 2105 2660 2109 2664
rect 2125 2660 2129 2664
rect 2185 2660 2189 2664
rect 2205 2660 2209 2664
rect 2265 2660 2269 2664
rect 2285 2660 2289 2664
rect 2331 2660 2335 2664
rect 2405 2660 2409 2664
rect 2425 2660 2429 2664
rect 2471 2660 2475 2664
rect 2531 2660 2535 2664
rect 2541 2660 2545 2664
rect 2561 2660 2565 2664
rect 2631 2660 2635 2664
rect 2651 2660 2655 2664
rect 2671 2660 2675 2664
rect 2731 2660 2735 2664
rect 2751 2660 2755 2664
rect 2771 2660 2775 2664
rect 2833 2660 2837 2664
rect 2843 2660 2847 2664
rect 2915 2660 2919 2664
rect 2935 2660 2939 2664
rect 2945 2660 2949 2664
rect 2967 2660 2971 2664
rect 2977 2660 2981 2664
rect 2999 2660 3003 2664
rect 3045 2660 3049 2664
rect 3053 2660 3057 2664
rect 3073 2660 3077 2664
rect 3083 2660 3087 2664
rect 3105 2660 3109 2664
rect 3155 2660 3159 2664
rect 3175 2660 3179 2664
rect 3185 2660 3189 2664
rect 3207 2660 3211 2664
rect 3217 2660 3221 2664
rect 3239 2660 3243 2664
rect 3285 2660 3289 2664
rect 3293 2660 3297 2664
rect 3313 2660 3317 2664
rect 3323 2660 3327 2664
rect 3345 2660 3349 2664
rect 3405 2660 3409 2664
rect 3465 2660 3469 2664
rect 3485 2660 3489 2664
rect 3545 2660 3549 2664
rect 3595 2660 3599 2664
rect 3615 2660 3619 2664
rect 3625 2660 3629 2664
rect 3647 2660 3651 2664
rect 3657 2660 3661 2664
rect 3679 2660 3683 2664
rect 3725 2660 3729 2664
rect 3733 2660 3737 2664
rect 3753 2660 3757 2664
rect 3763 2660 3767 2664
rect 3785 2660 3789 2664
rect 3866 2660 3870 2664
rect 3874 2660 3878 2664
rect 3894 2660 3898 2664
rect 3902 2660 3906 2664
rect 3965 2660 3969 2664
rect 3985 2660 3989 2664
rect 4031 2660 4035 2664
rect 4051 2660 4055 2664
rect 4071 2660 4075 2664
rect 4145 2660 4149 2664
rect 4165 2660 4169 2664
rect 4185 2660 4189 2664
rect 4231 2660 4235 2664
rect 4251 2660 4255 2664
rect 4315 2660 4319 2664
rect 4335 2660 4339 2664
rect 4345 2660 4349 2664
rect 4367 2660 4371 2664
rect 4377 2660 4381 2664
rect 4399 2660 4403 2664
rect 4445 2660 4449 2664
rect 4453 2660 4457 2664
rect 4473 2660 4477 2664
rect 4483 2660 4487 2664
rect 4505 2660 4509 2664
rect 4551 2660 4555 2664
rect 4571 2660 4575 2664
rect 4591 2660 4595 2664
rect 4653 2660 4657 2664
rect 4663 2660 4667 2664
rect 32 2636 36 2640
rect 40 2636 44 2640
rect 48 2636 52 2640
rect 134 2636 138 2640
rect 142 2636 146 2640
rect 164 2636 168 2640
rect 245 2636 249 2640
rect 315 2636 319 2640
rect 335 2636 339 2640
rect 345 2636 349 2640
rect 412 2636 416 2640
rect 434 2636 438 2640
rect 442 2636 446 2640
rect 528 2636 532 2640
rect 536 2636 540 2640
rect 544 2636 548 2640
rect 605 2636 609 2640
rect 625 2636 629 2640
rect 645 2636 649 2640
rect 705 2636 709 2640
rect 773 2636 777 2640
rect 783 2636 787 2640
rect 868 2636 872 2640
rect 876 2636 880 2640
rect 884 2636 888 2640
rect 945 2636 949 2640
rect 965 2636 969 2640
rect 985 2636 989 2640
rect 1033 2636 1037 2640
rect 1043 2636 1047 2640
rect 1148 2636 1152 2640
rect 1156 2636 1160 2640
rect 1164 2636 1168 2640
rect 1225 2636 1229 2640
rect 1285 2636 1289 2640
rect 1305 2636 1309 2640
rect 1325 2636 1329 2640
rect 1373 2636 1377 2640
rect 1383 2636 1387 2640
rect 1451 2636 1455 2640
rect 1533 2636 1537 2640
rect 1543 2636 1547 2640
rect 1595 2636 1599 2640
rect 1615 2636 1619 2640
rect 1625 2636 1629 2640
rect 1647 2636 1651 2640
rect 1657 2636 1661 2640
rect 1679 2636 1683 2640
rect 1725 2636 1729 2640
rect 1733 2636 1737 2640
rect 1753 2636 1757 2640
rect 1763 2636 1767 2640
rect 1785 2636 1789 2640
rect 1833 2636 1837 2640
rect 1843 2636 1847 2640
rect 1913 2636 1917 2640
rect 1923 2636 1927 2640
rect 1992 2636 1996 2640
rect 2000 2636 2004 2640
rect 2008 2636 2012 2640
rect 2091 2636 2095 2640
rect 2111 2636 2115 2640
rect 2185 2636 2189 2640
rect 2245 2636 2249 2640
rect 2265 2636 2269 2640
rect 2325 2636 2329 2640
rect 2385 2636 2389 2640
rect 2405 2636 2409 2640
rect 2425 2636 2429 2640
rect 2471 2636 2475 2640
rect 2491 2636 2495 2640
rect 2551 2636 2555 2640
rect 2561 2636 2565 2640
rect 2581 2636 2585 2640
rect 2651 2636 2655 2640
rect 2671 2636 2675 2640
rect 2691 2636 2695 2640
rect 2773 2636 2777 2640
rect 2783 2636 2787 2640
rect 2831 2636 2835 2640
rect 2851 2636 2855 2640
rect 2871 2636 2875 2640
rect 2933 2636 2937 2640
rect 2943 2636 2947 2640
rect 3011 2636 3015 2640
rect 3033 2636 3037 2640
rect 3091 2636 3095 2640
rect 3111 2636 3115 2640
rect 3131 2636 3135 2640
rect 3203 2636 3207 2640
rect 3225 2636 3229 2640
rect 3293 2636 3297 2640
rect 3303 2636 3307 2640
rect 3354 2636 3358 2640
rect 3362 2636 3366 2640
rect 3382 2636 3386 2640
rect 3390 2636 3394 2640
rect 3471 2636 3475 2640
rect 3493 2636 3497 2640
rect 3563 2636 3567 2640
rect 3585 2636 3589 2640
rect 3635 2636 3639 2640
rect 3655 2636 3659 2640
rect 3665 2636 3669 2640
rect 3687 2636 3691 2640
rect 3697 2636 3701 2640
rect 3719 2636 3723 2640
rect 3765 2636 3769 2640
rect 3773 2636 3777 2640
rect 3793 2636 3797 2640
rect 3803 2636 3807 2640
rect 3825 2636 3829 2640
rect 3892 2636 3896 2640
rect 3914 2636 3918 2640
rect 3922 2636 3926 2640
rect 3971 2636 3975 2640
rect 3991 2636 3995 2640
rect 4051 2636 4055 2640
rect 4071 2636 4075 2640
rect 4091 2636 4095 2640
rect 4111 2636 4115 2640
rect 4131 2636 4135 2640
rect 4151 2636 4155 2640
rect 4171 2636 4175 2640
rect 4191 2636 4195 2640
rect 4255 2636 4259 2640
rect 4275 2636 4279 2640
rect 4285 2636 4289 2640
rect 4307 2636 4311 2640
rect 4317 2636 4321 2640
rect 4339 2636 4343 2640
rect 4385 2636 4389 2640
rect 4393 2636 4397 2640
rect 4413 2636 4417 2640
rect 4423 2636 4427 2640
rect 4445 2636 4449 2640
rect 4491 2636 4495 2640
rect 4511 2636 4515 2640
rect 4531 2636 4535 2640
rect 4593 2636 4597 2640
rect 4603 2636 4607 2640
rect 4673 2636 4677 2640
rect 4683 2636 4687 2640
rect 134 2592 138 2596
rect 119 2586 138 2592
rect 32 2519 36 2576
rect 26 2507 36 2519
rect 20 2476 26 2507
rect 40 2499 44 2576
rect 48 2519 52 2576
rect 119 2573 126 2586
rect 119 2524 126 2561
rect 142 2559 146 2596
rect 164 2573 168 2616
rect 166 2561 175 2573
rect 140 2524 146 2547
rect 48 2507 55 2519
rect 67 2507 75 2519
rect 119 2518 135 2524
rect 140 2518 155 2524
rect 40 2480 46 2487
rect 40 2476 55 2480
rect 20 2472 35 2476
rect 31 2464 35 2472
rect 51 2464 55 2476
rect 71 2464 75 2507
rect 131 2504 135 2518
rect 151 2504 155 2518
rect 171 2504 175 2561
rect 245 2559 249 2616
rect 315 2590 319 2596
rect 301 2578 313 2590
rect 245 2547 254 2559
rect 245 2464 249 2547
rect 301 2504 305 2578
rect 335 2553 339 2596
rect 326 2541 339 2553
rect 323 2464 327 2541
rect 345 2539 349 2596
rect 412 2573 416 2616
rect 405 2561 414 2573
rect 345 2527 354 2539
rect 345 2464 349 2527
rect 405 2504 409 2561
rect 434 2559 438 2596
rect 442 2592 446 2596
rect 442 2586 461 2592
rect 454 2573 461 2586
rect 434 2524 440 2547
rect 454 2524 461 2561
rect 425 2518 440 2524
rect 445 2518 461 2524
rect 528 2519 532 2576
rect 425 2504 429 2518
rect 445 2504 449 2518
rect 505 2507 513 2519
rect 525 2507 532 2519
rect 505 2464 509 2507
rect 536 2499 540 2576
rect 544 2519 548 2576
rect 605 2519 609 2596
rect 625 2573 629 2596
rect 645 2591 649 2596
rect 645 2584 658 2591
rect 625 2561 634 2573
rect 544 2507 554 2519
rect 607 2507 614 2519
rect 534 2480 540 2487
rect 525 2476 540 2480
rect 554 2476 560 2507
rect 525 2464 529 2476
rect 545 2472 560 2476
rect 545 2464 549 2472
rect 610 2464 614 2507
rect 632 2504 636 2561
rect 654 2539 658 2584
rect 705 2573 709 2596
rect 773 2576 777 2596
rect 705 2561 714 2573
rect 763 2569 777 2576
rect 783 2576 787 2596
rect 783 2569 791 2576
rect 654 2516 658 2527
rect 640 2508 658 2516
rect 640 2504 644 2508
rect 705 2504 709 2561
rect 763 2553 769 2569
rect 766 2541 769 2553
rect 765 2464 769 2541
rect 785 2553 791 2569
rect 785 2541 794 2553
rect 785 2464 789 2541
rect 868 2519 872 2576
rect 845 2507 853 2519
rect 865 2507 872 2519
rect 845 2464 849 2507
rect 876 2499 880 2576
rect 884 2519 888 2576
rect 945 2519 949 2596
rect 965 2573 969 2596
rect 985 2591 989 2596
rect 985 2584 998 2591
rect 965 2561 974 2573
rect 884 2507 894 2519
rect 947 2507 954 2519
rect 874 2480 880 2487
rect 865 2476 880 2480
rect 894 2476 900 2507
rect 865 2464 869 2476
rect 885 2472 900 2476
rect 885 2464 889 2472
rect 950 2464 954 2507
rect 972 2504 976 2561
rect 994 2539 998 2584
rect 1033 2576 1037 2596
rect 1029 2569 1037 2576
rect 1043 2576 1047 2596
rect 1043 2569 1057 2576
rect 1029 2553 1035 2569
rect 1026 2541 1035 2553
rect 994 2516 998 2527
rect 980 2508 998 2516
rect 980 2504 984 2508
rect 1031 2464 1035 2541
rect 1051 2553 1057 2569
rect 1051 2541 1054 2553
rect 1051 2464 1055 2541
rect 1148 2519 1152 2576
rect 1125 2507 1133 2519
rect 1145 2507 1152 2519
rect 1125 2464 1129 2507
rect 1156 2499 1160 2576
rect 1164 2519 1168 2576
rect 1225 2559 1229 2616
rect 1225 2547 1234 2559
rect 1164 2507 1174 2519
rect 1154 2480 1160 2487
rect 1145 2476 1160 2480
rect 1174 2476 1180 2507
rect 1145 2464 1149 2476
rect 1165 2472 1180 2476
rect 1165 2464 1169 2472
rect 1225 2464 1229 2547
rect 1285 2519 1289 2596
rect 1305 2573 1309 2596
rect 1325 2591 1329 2596
rect 1325 2584 1338 2591
rect 1305 2561 1314 2573
rect 1287 2507 1294 2519
rect 1290 2464 1294 2507
rect 1312 2504 1316 2561
rect 1334 2539 1338 2584
rect 1373 2576 1377 2596
rect 1369 2569 1377 2576
rect 1383 2576 1387 2596
rect 1383 2569 1397 2576
rect 1451 2573 1455 2596
rect 1533 2576 1537 2596
rect 1369 2553 1375 2569
rect 1366 2541 1375 2553
rect 1334 2516 1338 2527
rect 1320 2508 1338 2516
rect 1320 2504 1324 2508
rect 1371 2464 1375 2541
rect 1391 2553 1397 2569
rect 1446 2561 1455 2573
rect 1391 2541 1394 2553
rect 1391 2464 1395 2541
rect 1451 2504 1455 2561
rect 1523 2569 1537 2576
rect 1543 2576 1547 2596
rect 1543 2569 1551 2576
rect 1523 2553 1529 2569
rect 1526 2541 1529 2553
rect 1525 2464 1529 2541
rect 1545 2553 1551 2569
rect 1595 2559 1599 2596
rect 1545 2541 1554 2553
rect 1615 2558 1619 2616
rect 1625 2584 1629 2616
rect 1647 2604 1651 2616
rect 1649 2592 1651 2604
rect 1657 2604 1661 2616
rect 1657 2592 1659 2604
rect 1625 2580 1658 2584
rect 1545 2464 1549 2541
rect 1595 2504 1599 2547
rect 1615 2464 1619 2546
rect 1634 2531 1638 2560
rect 1629 2523 1638 2531
rect 1629 2464 1633 2523
rect 1654 2516 1658 2580
rect 1655 2504 1658 2516
rect 1649 2464 1653 2504
rect 1663 2482 1667 2592
rect 1679 2502 1683 2616
rect 1725 2612 1729 2616
rect 1695 2608 1729 2612
rect 1661 2464 1665 2470
rect 1681 2464 1685 2490
rect 1695 2482 1699 2608
rect 1733 2604 1737 2616
rect 1707 2600 1737 2604
rect 1719 2599 1737 2600
rect 1753 2595 1757 2616
rect 1733 2591 1757 2595
rect 1733 2496 1739 2591
rect 1763 2567 1767 2616
rect 1763 2509 1767 2555
rect 1785 2528 1789 2596
rect 1833 2576 1837 2596
rect 1829 2569 1837 2576
rect 1843 2576 1847 2596
rect 1913 2576 1917 2596
rect 1843 2569 1857 2576
rect 1829 2553 1835 2569
rect 1826 2541 1835 2553
rect 1787 2516 1789 2528
rect 1763 2503 1771 2509
rect 1785 2504 1789 2516
rect 1707 2470 1731 2472
rect 1695 2468 1731 2470
rect 1727 2464 1731 2468
rect 1735 2464 1739 2496
rect 1755 2444 1759 2484
rect 1767 2474 1771 2503
rect 1763 2467 1771 2474
rect 1763 2444 1767 2467
rect 1831 2464 1835 2541
rect 1851 2553 1857 2569
rect 1909 2569 1917 2576
rect 1923 2576 1927 2596
rect 1923 2569 1937 2576
rect 1909 2553 1915 2569
rect 1851 2541 1854 2553
rect 1906 2541 1915 2553
rect 1851 2464 1855 2541
rect 1911 2464 1915 2541
rect 1931 2553 1937 2569
rect 1931 2541 1934 2553
rect 1931 2464 1935 2541
rect 1992 2519 1996 2576
rect 1986 2507 1996 2519
rect 1980 2476 1986 2507
rect 2000 2499 2004 2576
rect 2008 2519 2012 2576
rect 2091 2539 2095 2616
rect 2111 2539 2115 2616
rect 2185 2559 2189 2616
rect 2185 2547 2194 2559
rect 2086 2527 2095 2539
rect 2008 2507 2015 2519
rect 2027 2507 2035 2519
rect 2000 2480 2006 2487
rect 2000 2476 2015 2480
rect 1980 2472 1995 2476
rect 1991 2464 1995 2472
rect 2011 2464 2015 2476
rect 2031 2464 2035 2507
rect 2091 2504 2095 2527
rect 2099 2527 2114 2539
rect 2099 2504 2103 2527
rect 2185 2464 2189 2547
rect 2245 2539 2249 2616
rect 2265 2539 2269 2616
rect 2325 2559 2329 2616
rect 2325 2547 2334 2559
rect 2246 2527 2261 2539
rect 2257 2504 2261 2527
rect 2265 2527 2274 2539
rect 2265 2504 2269 2527
rect 2325 2464 2329 2547
rect 2385 2519 2389 2596
rect 2405 2573 2409 2596
rect 2425 2591 2429 2596
rect 2425 2584 2438 2591
rect 2405 2561 2414 2573
rect 2387 2507 2394 2519
rect 2390 2464 2394 2507
rect 2412 2504 2416 2561
rect 2434 2539 2438 2584
rect 2471 2539 2475 2616
rect 2491 2539 2495 2616
rect 2831 2609 2835 2616
rect 2851 2609 2855 2616
rect 2822 2604 2835 2609
rect 2551 2539 2555 2596
rect 2561 2553 2565 2596
rect 2581 2590 2585 2596
rect 2651 2591 2655 2596
rect 2587 2578 2599 2590
rect 2561 2541 2574 2553
rect 2466 2527 2475 2539
rect 2434 2516 2438 2527
rect 2420 2508 2438 2516
rect 2420 2504 2424 2508
rect 2471 2504 2475 2527
rect 2479 2527 2494 2539
rect 2546 2527 2555 2539
rect 2479 2504 2483 2527
rect 2551 2464 2555 2527
rect 2573 2464 2577 2541
rect 2595 2504 2599 2578
rect 2642 2584 2655 2591
rect 2642 2539 2646 2584
rect 2671 2573 2675 2596
rect 2666 2561 2675 2573
rect 2642 2516 2646 2527
rect 2642 2508 2660 2516
rect 2656 2504 2660 2508
rect 2664 2504 2668 2561
rect 2691 2519 2695 2596
rect 2773 2576 2777 2596
rect 2763 2569 2777 2576
rect 2783 2576 2787 2596
rect 2783 2569 2791 2576
rect 2763 2553 2769 2569
rect 2766 2541 2769 2553
rect 2686 2507 2693 2519
rect 2686 2464 2690 2507
rect 2765 2464 2769 2541
rect 2785 2553 2791 2569
rect 2822 2559 2826 2604
rect 2785 2541 2794 2553
rect 2785 2464 2789 2541
rect 2822 2513 2826 2547
rect 2841 2603 2855 2609
rect 2841 2539 2845 2603
rect 2871 2588 2875 2596
rect 2865 2576 2875 2588
rect 2933 2576 2937 2596
rect 2929 2569 2937 2576
rect 2943 2576 2947 2596
rect 2943 2569 2957 2576
rect 2929 2553 2935 2569
rect 2926 2541 2935 2553
rect 2822 2508 2835 2513
rect 2831 2504 2835 2508
rect 2841 2504 2845 2527
rect 2861 2504 2865 2509
rect 2931 2464 2935 2541
rect 2951 2553 2957 2569
rect 2951 2541 2954 2553
rect 2951 2464 2955 2541
rect 3011 2539 3015 2616
rect 3033 2590 3037 2596
rect 3091 2591 3095 2596
rect 3035 2578 3037 2590
rect 3082 2584 3095 2591
rect 3082 2539 3086 2584
rect 3111 2573 3115 2596
rect 3106 2561 3115 2573
rect 3006 2527 3015 2539
rect 3011 2464 3015 2527
rect 3035 2510 3037 2522
rect 3033 2504 3037 2510
rect 3082 2516 3086 2527
rect 3082 2508 3100 2516
rect 3096 2504 3100 2508
rect 3104 2504 3108 2561
rect 3131 2519 3135 2596
rect 3203 2590 3207 2596
rect 3203 2578 3205 2590
rect 3225 2539 3229 2616
rect 3293 2576 3297 2596
rect 3283 2569 3297 2576
rect 3303 2576 3307 2596
rect 3354 2588 3358 2596
rect 3341 2581 3358 2588
rect 3303 2569 3311 2576
rect 3283 2553 3289 2569
rect 3286 2541 3289 2553
rect 3225 2527 3234 2539
rect 3126 2507 3133 2519
rect 3203 2510 3205 2522
rect 3126 2464 3130 2507
rect 3203 2504 3207 2510
rect 3225 2464 3229 2527
rect 3285 2464 3289 2541
rect 3305 2553 3311 2569
rect 3305 2541 3314 2553
rect 3305 2464 3309 2541
rect 3341 2539 3347 2581
rect 3362 2573 3366 2596
rect 3382 2582 3386 2596
rect 3390 2591 3394 2596
rect 3390 2587 3420 2591
rect 3382 2575 3395 2582
rect 3391 2573 3395 2575
rect 3391 2561 3393 2573
rect 3362 2532 3366 2561
rect 3347 2527 3355 2532
rect 3335 2526 3355 2527
rect 3362 2526 3375 2532
rect 3351 2504 3355 2526
rect 3371 2504 3375 2526
rect 3391 2504 3395 2561
rect 3414 2539 3420 2587
rect 3471 2539 3475 2616
rect 3493 2590 3497 2596
rect 3495 2578 3497 2590
rect 3563 2590 3567 2596
rect 3563 2578 3565 2590
rect 3411 2527 3414 2539
rect 3466 2527 3475 2539
rect 3411 2504 3415 2527
rect 3471 2464 3475 2527
rect 3585 2539 3589 2616
rect 3635 2559 3639 2596
rect 3655 2558 3659 2616
rect 3665 2584 3669 2616
rect 3687 2604 3691 2616
rect 3689 2592 3691 2604
rect 3697 2604 3701 2616
rect 3697 2592 3699 2604
rect 3665 2580 3698 2584
rect 3585 2527 3594 2539
rect 3495 2510 3497 2522
rect 3493 2504 3497 2510
rect 3563 2510 3565 2522
rect 3563 2504 3567 2510
rect 3585 2464 3589 2527
rect 3635 2504 3639 2547
rect 3655 2464 3659 2546
rect 3674 2531 3678 2560
rect 3669 2523 3678 2531
rect 3669 2464 3673 2523
rect 3694 2516 3698 2580
rect 3695 2504 3698 2516
rect 3689 2464 3693 2504
rect 3703 2482 3707 2592
rect 3719 2502 3723 2616
rect 3765 2612 3769 2616
rect 3735 2608 3769 2612
rect 3701 2464 3705 2470
rect 3721 2464 3725 2490
rect 3735 2482 3739 2608
rect 3773 2604 3777 2616
rect 3747 2600 3777 2604
rect 3759 2599 3777 2600
rect 3793 2595 3797 2616
rect 3773 2591 3797 2595
rect 3773 2496 3779 2591
rect 3803 2567 3807 2616
rect 3803 2509 3807 2555
rect 3825 2528 3829 2596
rect 3892 2573 3896 2616
rect 3827 2516 3829 2528
rect 3803 2503 3811 2509
rect 3825 2504 3829 2516
rect 3885 2561 3894 2573
rect 3885 2504 3889 2561
rect 3914 2559 3918 2596
rect 3922 2592 3926 2596
rect 3922 2586 3941 2592
rect 3934 2573 3941 2586
rect 3914 2524 3920 2547
rect 3934 2524 3941 2561
rect 3971 2539 3975 2616
rect 3991 2539 3995 2616
rect 4051 2573 4055 2596
rect 4071 2573 4075 2596
rect 4091 2576 4095 2596
rect 4111 2576 4115 2596
rect 4131 2576 4135 2596
rect 4151 2576 4155 2596
rect 4171 2576 4175 2596
rect 4191 2576 4195 2596
rect 4051 2561 4054 2573
rect 4066 2561 4075 2573
rect 4102 2564 4115 2576
rect 4142 2564 4155 2576
rect 4182 2564 4195 2576
rect 3966 2527 3975 2539
rect 3905 2518 3920 2524
rect 3925 2518 3941 2524
rect 3905 2504 3909 2518
rect 3925 2504 3929 2518
rect 3971 2504 3975 2527
rect 3979 2527 3994 2539
rect 3979 2504 3983 2527
rect 4051 2504 4055 2561
rect 4071 2504 4075 2561
rect 4091 2504 4095 2564
rect 4111 2504 4115 2564
rect 4131 2504 4135 2564
rect 4151 2504 4155 2564
rect 4171 2504 4175 2564
rect 4191 2504 4195 2564
rect 4255 2559 4259 2596
rect 4275 2558 4279 2616
rect 4285 2584 4289 2616
rect 4307 2604 4311 2616
rect 4309 2592 4311 2604
rect 4317 2604 4321 2616
rect 4317 2592 4319 2604
rect 4285 2580 4318 2584
rect 4255 2504 4259 2547
rect 3747 2470 3771 2472
rect 3735 2468 3771 2470
rect 3767 2464 3771 2468
rect 3775 2464 3779 2496
rect 3795 2444 3799 2484
rect 3807 2474 3811 2503
rect 3803 2467 3811 2474
rect 3803 2444 3807 2467
rect 4275 2464 4279 2546
rect 4294 2531 4298 2560
rect 4289 2523 4298 2531
rect 4289 2464 4293 2523
rect 4314 2516 4318 2580
rect 4315 2504 4318 2516
rect 4309 2464 4313 2504
rect 4323 2482 4327 2592
rect 4339 2502 4343 2616
rect 4385 2612 4389 2616
rect 4355 2608 4389 2612
rect 4321 2464 4325 2470
rect 4341 2464 4345 2490
rect 4355 2482 4359 2608
rect 4393 2604 4397 2616
rect 4367 2600 4397 2604
rect 4379 2599 4397 2600
rect 4413 2595 4417 2616
rect 4393 2591 4417 2595
rect 4393 2496 4399 2591
rect 4423 2567 4427 2616
rect 4423 2509 4427 2555
rect 4445 2528 4449 2596
rect 4491 2591 4495 2596
rect 4482 2584 4495 2591
rect 4482 2539 4486 2584
rect 4511 2573 4515 2596
rect 4506 2561 4515 2573
rect 4447 2516 4449 2528
rect 4423 2503 4431 2509
rect 4445 2504 4449 2516
rect 4482 2516 4486 2527
rect 4482 2508 4500 2516
rect 4496 2504 4500 2508
rect 4504 2504 4508 2561
rect 4531 2519 4535 2596
rect 4593 2576 4597 2596
rect 4589 2569 4597 2576
rect 4603 2576 4607 2596
rect 4673 2576 4677 2596
rect 4603 2569 4617 2576
rect 4589 2553 4595 2569
rect 4586 2541 4595 2553
rect 4526 2507 4533 2519
rect 4367 2470 4391 2472
rect 4355 2468 4391 2470
rect 4387 2464 4391 2468
rect 4395 2464 4399 2496
rect 4415 2444 4419 2484
rect 4427 2474 4431 2503
rect 4423 2467 4431 2474
rect 4423 2444 4427 2467
rect 4526 2464 4530 2507
rect 4591 2464 4595 2541
rect 4611 2553 4617 2569
rect 4669 2569 4677 2576
rect 4683 2576 4687 2596
rect 4683 2569 4697 2576
rect 4669 2553 4675 2569
rect 4611 2541 4614 2553
rect 4666 2541 4675 2553
rect 4611 2464 4615 2541
rect 4671 2464 4675 2541
rect 4691 2553 4697 2569
rect 4691 2541 4694 2553
rect 4691 2464 4695 2541
rect 31 2420 35 2424
rect 51 2420 55 2424
rect 71 2420 75 2424
rect 131 2420 135 2424
rect 151 2420 155 2424
rect 171 2420 175 2424
rect 245 2420 249 2424
rect 301 2420 305 2424
rect 323 2420 327 2424
rect 345 2420 349 2424
rect 405 2420 409 2424
rect 425 2420 429 2424
rect 445 2420 449 2424
rect 505 2420 509 2424
rect 525 2420 529 2424
rect 545 2420 549 2424
rect 610 2420 614 2424
rect 632 2420 636 2424
rect 640 2420 644 2424
rect 705 2420 709 2424
rect 765 2420 769 2424
rect 785 2420 789 2424
rect 845 2420 849 2424
rect 865 2420 869 2424
rect 885 2420 889 2424
rect 950 2420 954 2424
rect 972 2420 976 2424
rect 980 2420 984 2424
rect 1031 2420 1035 2424
rect 1051 2420 1055 2424
rect 1125 2420 1129 2424
rect 1145 2420 1149 2424
rect 1165 2420 1169 2424
rect 1225 2420 1229 2424
rect 1290 2420 1294 2424
rect 1312 2420 1316 2424
rect 1320 2420 1324 2424
rect 1371 2420 1375 2424
rect 1391 2420 1395 2424
rect 1451 2420 1455 2424
rect 1525 2420 1529 2424
rect 1545 2420 1549 2424
rect 1595 2420 1599 2424
rect 1615 2420 1619 2424
rect 1629 2420 1633 2424
rect 1649 2420 1653 2424
rect 1661 2420 1665 2424
rect 1681 2420 1685 2424
rect 1727 2420 1731 2424
rect 1735 2420 1739 2424
rect 1755 2420 1759 2424
rect 1763 2420 1767 2424
rect 1785 2420 1789 2424
rect 1831 2420 1835 2424
rect 1851 2420 1855 2424
rect 1911 2420 1915 2424
rect 1931 2420 1935 2424
rect 1991 2420 1995 2424
rect 2011 2420 2015 2424
rect 2031 2420 2035 2424
rect 2091 2420 2095 2424
rect 2099 2420 2103 2424
rect 2185 2420 2189 2424
rect 2257 2420 2261 2424
rect 2265 2420 2269 2424
rect 2325 2420 2329 2424
rect 2390 2420 2394 2424
rect 2412 2420 2416 2424
rect 2420 2420 2424 2424
rect 2471 2420 2475 2424
rect 2479 2420 2483 2424
rect 2551 2420 2555 2424
rect 2573 2420 2577 2424
rect 2595 2420 2599 2424
rect 2656 2420 2660 2424
rect 2664 2420 2668 2424
rect 2686 2420 2690 2424
rect 2765 2420 2769 2424
rect 2785 2420 2789 2424
rect 2831 2420 2835 2424
rect 2841 2420 2845 2424
rect 2861 2420 2865 2424
rect 2931 2420 2935 2424
rect 2951 2420 2955 2424
rect 3011 2420 3015 2424
rect 3033 2420 3037 2424
rect 3096 2420 3100 2424
rect 3104 2420 3108 2424
rect 3126 2420 3130 2424
rect 3203 2420 3207 2424
rect 3225 2420 3229 2424
rect 3285 2420 3289 2424
rect 3305 2420 3309 2424
rect 3351 2420 3355 2424
rect 3371 2420 3375 2424
rect 3391 2420 3395 2424
rect 3411 2420 3415 2424
rect 3471 2420 3475 2424
rect 3493 2420 3497 2424
rect 3563 2420 3567 2424
rect 3585 2420 3589 2424
rect 3635 2420 3639 2424
rect 3655 2420 3659 2424
rect 3669 2420 3673 2424
rect 3689 2420 3693 2424
rect 3701 2420 3705 2424
rect 3721 2420 3725 2424
rect 3767 2420 3771 2424
rect 3775 2420 3779 2424
rect 3795 2420 3799 2424
rect 3803 2420 3807 2424
rect 3825 2420 3829 2424
rect 3885 2420 3889 2424
rect 3905 2420 3909 2424
rect 3925 2420 3929 2424
rect 3971 2420 3975 2424
rect 3979 2420 3983 2424
rect 4051 2420 4055 2424
rect 4071 2420 4075 2424
rect 4091 2420 4095 2424
rect 4111 2420 4115 2424
rect 4131 2420 4135 2424
rect 4151 2420 4155 2424
rect 4171 2420 4175 2424
rect 4191 2420 4195 2424
rect 4255 2420 4259 2424
rect 4275 2420 4279 2424
rect 4289 2420 4293 2424
rect 4309 2420 4313 2424
rect 4321 2420 4325 2424
rect 4341 2420 4345 2424
rect 4387 2420 4391 2424
rect 4395 2420 4399 2424
rect 4415 2420 4419 2424
rect 4423 2420 4427 2424
rect 4445 2420 4449 2424
rect 4496 2420 4500 2424
rect 4504 2420 4508 2424
rect 4526 2420 4530 2424
rect 4591 2420 4595 2424
rect 4611 2420 4615 2424
rect 4671 2420 4675 2424
rect 4691 2420 4695 2424
rect 45 2396 49 2400
rect 65 2396 69 2400
rect 85 2396 89 2400
rect 150 2396 154 2400
rect 172 2396 176 2400
rect 180 2396 184 2400
rect 236 2396 240 2400
rect 244 2396 248 2400
rect 266 2396 270 2400
rect 331 2396 335 2400
rect 351 2396 355 2400
rect 371 2396 375 2400
rect 431 2396 435 2400
rect 451 2396 455 2400
rect 471 2396 475 2400
rect 536 2396 540 2400
rect 544 2396 548 2400
rect 566 2396 570 2400
rect 645 2396 649 2400
rect 665 2396 669 2400
rect 685 2396 689 2400
rect 731 2396 735 2400
rect 801 2396 805 2400
rect 823 2396 827 2400
rect 845 2396 849 2400
rect 891 2396 895 2400
rect 911 2396 915 2400
rect 971 2396 975 2400
rect 993 2396 997 2400
rect 1015 2396 1019 2400
rect 1090 2396 1094 2400
rect 1112 2396 1116 2400
rect 1120 2396 1124 2400
rect 1190 2396 1194 2400
rect 1212 2396 1216 2400
rect 1220 2396 1224 2400
rect 1275 2396 1279 2400
rect 1295 2396 1299 2400
rect 1309 2396 1313 2400
rect 1329 2396 1333 2400
rect 1341 2396 1345 2400
rect 1361 2396 1365 2400
rect 1407 2396 1411 2400
rect 1415 2396 1419 2400
rect 1435 2396 1439 2400
rect 1443 2396 1447 2400
rect 1465 2396 1469 2400
rect 1530 2396 1534 2400
rect 1552 2396 1556 2400
rect 1560 2396 1564 2400
rect 1615 2396 1619 2400
rect 1635 2396 1639 2400
rect 1649 2396 1653 2400
rect 1669 2396 1673 2400
rect 1681 2396 1685 2400
rect 1701 2396 1705 2400
rect 1747 2396 1751 2400
rect 1755 2396 1759 2400
rect 1775 2396 1779 2400
rect 1783 2396 1787 2400
rect 1805 2396 1809 2400
rect 1865 2396 1869 2400
rect 1925 2396 1929 2400
rect 1976 2396 1980 2400
rect 1984 2396 1988 2400
rect 2006 2396 2010 2400
rect 2075 2396 2079 2400
rect 2095 2396 2099 2400
rect 2109 2396 2113 2400
rect 2129 2396 2133 2400
rect 2141 2396 2145 2400
rect 2161 2396 2165 2400
rect 2207 2396 2211 2400
rect 2215 2396 2219 2400
rect 2235 2396 2239 2400
rect 2243 2396 2247 2400
rect 2265 2396 2269 2400
rect 2325 2396 2329 2400
rect 2345 2396 2349 2400
rect 2365 2396 2369 2400
rect 2425 2396 2429 2400
rect 2445 2396 2449 2400
rect 2465 2396 2469 2400
rect 2511 2396 2515 2400
rect 2531 2396 2535 2400
rect 2551 2396 2555 2400
rect 2611 2396 2615 2400
rect 2633 2396 2637 2400
rect 2655 2396 2659 2400
rect 2711 2396 2715 2400
rect 2733 2396 2737 2400
rect 2741 2396 2745 2400
rect 2761 2396 2765 2400
rect 2769 2396 2773 2400
rect 2815 2396 2819 2400
rect 2835 2396 2839 2400
rect 2847 2396 2851 2400
rect 2867 2396 2871 2400
rect 2881 2396 2885 2400
rect 2901 2396 2905 2400
rect 2970 2396 2974 2400
rect 2992 2396 2996 2400
rect 3000 2396 3004 2400
rect 3070 2396 3074 2400
rect 3092 2396 3096 2400
rect 3100 2396 3104 2400
rect 3156 2396 3160 2400
rect 3164 2396 3168 2400
rect 3186 2396 3190 2400
rect 3251 2396 3255 2400
rect 3273 2396 3277 2400
rect 3281 2396 3285 2400
rect 3301 2396 3305 2400
rect 3309 2396 3313 2400
rect 3355 2396 3359 2400
rect 3375 2396 3379 2400
rect 3387 2396 3391 2400
rect 3407 2396 3411 2400
rect 3421 2396 3425 2400
rect 3441 2396 3445 2400
rect 3510 2396 3514 2400
rect 3532 2396 3536 2400
rect 3540 2396 3544 2400
rect 3617 2396 3621 2400
rect 3625 2396 3629 2400
rect 3671 2396 3675 2400
rect 3681 2396 3685 2400
rect 3701 2396 3705 2400
rect 3785 2396 3789 2400
rect 3805 2396 3809 2400
rect 3865 2396 3869 2400
rect 3885 2396 3889 2400
rect 3905 2396 3909 2400
rect 3925 2396 3929 2400
rect 3985 2396 3989 2400
rect 4005 2396 4009 2400
rect 4025 2396 4029 2400
rect 4045 2396 4049 2400
rect 4095 2396 4099 2400
rect 4115 2396 4119 2400
rect 4129 2396 4133 2400
rect 4149 2396 4153 2400
rect 4161 2396 4165 2400
rect 4181 2396 4185 2400
rect 4227 2396 4231 2400
rect 4235 2396 4239 2400
rect 4255 2396 4259 2400
rect 4263 2396 4267 2400
rect 4285 2396 4289 2400
rect 4331 2396 4335 2400
rect 4353 2396 4357 2400
rect 4361 2396 4365 2400
rect 4381 2396 4385 2400
rect 4389 2396 4393 2400
rect 4435 2396 4439 2400
rect 4455 2396 4459 2400
rect 4467 2396 4471 2400
rect 4487 2396 4491 2400
rect 4501 2396 4505 2400
rect 4521 2396 4525 2400
rect 4576 2396 4580 2400
rect 4584 2396 4588 2400
rect 4606 2396 4610 2400
rect 4671 2396 4675 2400
rect 4691 2396 4695 2400
rect 45 2313 49 2356
rect 65 2344 69 2356
rect 85 2348 89 2356
rect 85 2344 100 2348
rect 65 2340 80 2344
rect 74 2333 80 2340
rect 45 2301 53 2313
rect 65 2301 72 2313
rect 68 2244 72 2301
rect 76 2244 80 2321
rect 94 2313 100 2344
rect 150 2313 154 2356
rect 84 2301 94 2313
rect 147 2301 154 2313
rect 84 2244 88 2301
rect 145 2224 149 2301
rect 172 2259 176 2316
rect 180 2312 184 2316
rect 236 2312 240 2316
rect 180 2304 198 2312
rect 194 2293 198 2304
rect 222 2304 240 2312
rect 222 2293 226 2304
rect 165 2247 174 2259
rect 165 2224 169 2247
rect 194 2236 198 2281
rect 185 2229 198 2236
rect 222 2236 226 2281
rect 244 2259 248 2316
rect 266 2313 270 2356
rect 331 2348 335 2356
rect 320 2344 335 2348
rect 351 2344 355 2356
rect 320 2313 326 2344
rect 340 2340 355 2344
rect 340 2333 346 2340
rect 266 2301 273 2313
rect 326 2301 336 2313
rect 246 2247 255 2259
rect 222 2229 235 2236
rect 185 2224 189 2229
rect 231 2224 235 2229
rect 251 2224 255 2247
rect 271 2224 275 2301
rect 332 2244 336 2301
rect 340 2244 344 2321
rect 371 2313 375 2356
rect 348 2301 355 2313
rect 367 2301 375 2313
rect 431 2302 435 2316
rect 451 2302 455 2316
rect 348 2244 352 2301
rect 419 2296 435 2302
rect 440 2296 455 2302
rect 419 2259 426 2296
rect 440 2273 446 2296
rect 419 2234 426 2247
rect 419 2228 438 2234
rect 434 2224 438 2228
rect 442 2224 446 2261
rect 471 2259 475 2316
rect 536 2312 540 2316
rect 522 2304 540 2312
rect 522 2293 526 2304
rect 466 2247 475 2259
rect 464 2204 468 2247
rect 522 2236 526 2281
rect 544 2259 548 2316
rect 566 2313 570 2356
rect 566 2301 573 2313
rect 546 2247 555 2259
rect 522 2229 535 2236
rect 531 2224 535 2229
rect 551 2224 555 2247
rect 571 2224 575 2301
rect 645 2259 649 2316
rect 665 2302 669 2316
rect 685 2302 689 2316
rect 665 2296 680 2302
rect 685 2296 701 2302
rect 674 2273 680 2296
rect 645 2247 654 2259
rect 652 2204 656 2247
rect 674 2224 678 2261
rect 694 2259 701 2296
rect 731 2273 735 2356
rect 726 2261 735 2273
rect 694 2234 701 2247
rect 682 2228 701 2234
rect 682 2224 686 2228
rect 731 2204 735 2261
rect 801 2242 805 2316
rect 823 2279 827 2356
rect 845 2293 849 2356
rect 845 2281 854 2293
rect 826 2267 839 2279
rect 801 2230 813 2242
rect 815 2224 819 2230
rect 835 2224 839 2267
rect 845 2224 849 2281
rect 891 2279 895 2356
rect 886 2267 895 2279
rect 889 2251 895 2267
rect 911 2279 915 2356
rect 971 2293 975 2356
rect 966 2281 975 2293
rect 911 2267 914 2279
rect 911 2251 917 2267
rect 889 2244 897 2251
rect 893 2224 897 2244
rect 903 2244 917 2251
rect 903 2224 907 2244
rect 971 2224 975 2281
rect 993 2279 997 2356
rect 981 2267 994 2279
rect 981 2224 985 2267
rect 1015 2242 1019 2316
rect 1090 2313 1094 2356
rect 1087 2301 1094 2313
rect 1007 2230 1019 2242
rect 1001 2224 1005 2230
rect 1085 2224 1089 2301
rect 1112 2259 1116 2316
rect 1120 2312 1124 2316
rect 1190 2313 1194 2356
rect 1120 2304 1138 2312
rect 1134 2293 1138 2304
rect 1187 2301 1194 2313
rect 1105 2247 1114 2259
rect 1105 2224 1109 2247
rect 1134 2236 1138 2281
rect 1125 2229 1138 2236
rect 1125 2224 1129 2229
rect 1185 2224 1189 2301
rect 1212 2259 1216 2316
rect 1220 2312 1224 2316
rect 1220 2304 1238 2312
rect 1234 2293 1238 2304
rect 1205 2247 1214 2259
rect 1205 2224 1209 2247
rect 1234 2236 1238 2281
rect 1275 2273 1279 2316
rect 1295 2274 1299 2356
rect 1309 2297 1313 2356
rect 1329 2316 1333 2356
rect 1341 2350 1345 2356
rect 1335 2304 1338 2316
rect 1309 2289 1318 2297
rect 1225 2229 1238 2236
rect 1225 2224 1229 2229
rect 1275 2224 1279 2261
rect 1295 2204 1299 2262
rect 1314 2260 1318 2289
rect 1334 2240 1338 2304
rect 1305 2236 1338 2240
rect 1305 2204 1309 2236
rect 1343 2228 1347 2338
rect 1361 2330 1365 2356
rect 1407 2352 1411 2356
rect 1375 2350 1411 2352
rect 1387 2348 1411 2350
rect 1329 2216 1331 2228
rect 1327 2204 1331 2216
rect 1337 2216 1339 2228
rect 1337 2204 1341 2216
rect 1359 2204 1363 2318
rect 1375 2212 1379 2338
rect 1415 2324 1419 2356
rect 1435 2336 1439 2376
rect 1443 2353 1447 2376
rect 1443 2346 1451 2353
rect 1413 2229 1419 2324
rect 1447 2317 1451 2346
rect 1443 2311 1451 2317
rect 1443 2265 1447 2311
rect 1465 2304 1469 2316
rect 1530 2313 1534 2356
rect 1467 2292 1469 2304
rect 1527 2301 1534 2313
rect 1413 2225 1437 2229
rect 1399 2220 1417 2221
rect 1387 2216 1417 2220
rect 1375 2208 1409 2212
rect 1405 2204 1409 2208
rect 1413 2204 1417 2216
rect 1433 2204 1437 2225
rect 1443 2204 1447 2253
rect 1465 2224 1469 2292
rect 1525 2224 1529 2301
rect 1552 2259 1556 2316
rect 1560 2312 1564 2316
rect 1560 2304 1578 2312
rect 1574 2293 1578 2304
rect 1545 2247 1554 2259
rect 1545 2224 1549 2247
rect 1574 2236 1578 2281
rect 1615 2273 1619 2316
rect 1635 2274 1639 2356
rect 1649 2297 1653 2356
rect 1669 2316 1673 2356
rect 1681 2350 1685 2356
rect 1675 2304 1678 2316
rect 1649 2289 1658 2297
rect 1565 2229 1578 2236
rect 1565 2224 1569 2229
rect 1615 2224 1619 2261
rect 1635 2204 1639 2262
rect 1654 2260 1658 2289
rect 1674 2240 1678 2304
rect 1645 2236 1678 2240
rect 1645 2204 1649 2236
rect 1683 2228 1687 2338
rect 1701 2330 1705 2356
rect 1747 2352 1751 2356
rect 1715 2350 1751 2352
rect 1727 2348 1751 2350
rect 1669 2216 1671 2228
rect 1667 2204 1671 2216
rect 1677 2216 1679 2228
rect 1677 2204 1681 2216
rect 1699 2204 1703 2318
rect 1715 2212 1719 2338
rect 1755 2324 1759 2356
rect 1775 2336 1779 2376
rect 1783 2353 1787 2376
rect 1783 2346 1791 2353
rect 1753 2229 1759 2324
rect 1787 2317 1791 2346
rect 1783 2311 1791 2317
rect 1783 2265 1787 2311
rect 1805 2304 1809 2316
rect 1807 2292 1809 2304
rect 1753 2225 1777 2229
rect 1739 2220 1757 2221
rect 1727 2216 1757 2220
rect 1715 2208 1749 2212
rect 1745 2204 1749 2208
rect 1753 2204 1757 2216
rect 1773 2204 1777 2225
rect 1783 2204 1787 2253
rect 1805 2224 1809 2292
rect 1865 2273 1869 2356
rect 1925 2273 1929 2356
rect 1976 2312 1980 2316
rect 1962 2304 1980 2312
rect 1962 2293 1966 2304
rect 1865 2261 1874 2273
rect 1925 2261 1934 2273
rect 1865 2204 1869 2261
rect 1925 2204 1929 2261
rect 1962 2236 1966 2281
rect 1984 2259 1988 2316
rect 2006 2313 2010 2356
rect 2006 2301 2013 2313
rect 1986 2247 1995 2259
rect 1962 2229 1975 2236
rect 1971 2224 1975 2229
rect 1991 2224 1995 2247
rect 2011 2224 2015 2301
rect 2075 2273 2079 2316
rect 2095 2274 2099 2356
rect 2109 2297 2113 2356
rect 2129 2316 2133 2356
rect 2141 2350 2145 2356
rect 2135 2304 2138 2316
rect 2109 2289 2118 2297
rect 2075 2224 2079 2261
rect 2095 2204 2099 2262
rect 2114 2260 2118 2289
rect 2134 2240 2138 2304
rect 2105 2236 2138 2240
rect 2105 2204 2109 2236
rect 2143 2228 2147 2338
rect 2161 2330 2165 2356
rect 2207 2352 2211 2356
rect 2175 2350 2211 2352
rect 2187 2348 2211 2350
rect 2129 2216 2131 2228
rect 2127 2204 2131 2216
rect 2137 2216 2139 2228
rect 2137 2204 2141 2216
rect 2159 2204 2163 2318
rect 2175 2212 2179 2338
rect 2215 2324 2219 2356
rect 2235 2336 2239 2376
rect 2243 2353 2247 2376
rect 2243 2346 2251 2353
rect 2213 2229 2219 2324
rect 2247 2317 2251 2346
rect 2243 2311 2251 2317
rect 2511 2348 2515 2356
rect 2500 2344 2515 2348
rect 2531 2344 2535 2356
rect 2243 2265 2247 2311
rect 2265 2304 2269 2316
rect 2267 2292 2269 2304
rect 2213 2225 2237 2229
rect 2199 2220 2217 2221
rect 2187 2216 2217 2220
rect 2175 2208 2209 2212
rect 2205 2204 2209 2208
rect 2213 2204 2217 2216
rect 2233 2204 2237 2225
rect 2243 2204 2247 2253
rect 2265 2224 2269 2292
rect 2325 2259 2329 2316
rect 2345 2302 2349 2316
rect 2365 2302 2369 2316
rect 2345 2296 2360 2302
rect 2365 2296 2381 2302
rect 2354 2273 2360 2296
rect 2325 2247 2334 2259
rect 2332 2204 2336 2247
rect 2354 2224 2358 2261
rect 2374 2259 2381 2296
rect 2425 2259 2429 2316
rect 2445 2302 2449 2316
rect 2465 2302 2469 2316
rect 2500 2313 2506 2344
rect 2520 2340 2535 2344
rect 2520 2333 2526 2340
rect 2445 2296 2460 2302
rect 2465 2296 2481 2302
rect 2506 2301 2516 2313
rect 2454 2273 2460 2296
rect 2425 2247 2434 2259
rect 2374 2234 2381 2247
rect 2362 2228 2381 2234
rect 2362 2224 2366 2228
rect 2432 2204 2436 2247
rect 2454 2224 2458 2261
rect 2474 2259 2481 2296
rect 2474 2234 2481 2247
rect 2512 2244 2516 2301
rect 2520 2244 2524 2321
rect 2551 2313 2555 2356
rect 2528 2301 2535 2313
rect 2547 2301 2555 2313
rect 2528 2244 2532 2301
rect 2611 2293 2615 2356
rect 2606 2281 2615 2293
rect 2462 2228 2481 2234
rect 2462 2224 2466 2228
rect 2611 2224 2615 2281
rect 2633 2279 2637 2356
rect 2733 2353 2737 2376
rect 2729 2346 2737 2353
rect 2729 2317 2733 2346
rect 2741 2336 2745 2376
rect 2761 2324 2765 2356
rect 2769 2352 2773 2356
rect 2769 2350 2805 2352
rect 2769 2348 2793 2350
rect 2621 2267 2634 2279
rect 2621 2224 2625 2267
rect 2655 2242 2659 2316
rect 2647 2230 2659 2242
rect 2711 2304 2715 2316
rect 2729 2311 2737 2317
rect 2711 2292 2713 2304
rect 2641 2224 2645 2230
rect 2711 2224 2715 2292
rect 2733 2265 2737 2311
rect 2733 2204 2737 2253
rect 2761 2229 2767 2324
rect 2743 2225 2767 2229
rect 2743 2204 2747 2225
rect 2763 2220 2781 2221
rect 2763 2216 2793 2220
rect 2763 2204 2767 2216
rect 2801 2212 2805 2338
rect 2815 2330 2819 2356
rect 2835 2350 2839 2356
rect 2771 2208 2805 2212
rect 2771 2204 2775 2208
rect 2817 2204 2821 2318
rect 2833 2228 2837 2338
rect 2847 2316 2851 2356
rect 2842 2304 2845 2316
rect 2842 2240 2846 2304
rect 2867 2297 2871 2356
rect 2862 2289 2871 2297
rect 2862 2260 2866 2289
rect 2881 2274 2885 2356
rect 2901 2273 2905 2316
rect 2970 2313 2974 2356
rect 2967 2301 2974 2313
rect 2842 2236 2875 2240
rect 2841 2216 2843 2228
rect 2839 2204 2843 2216
rect 2849 2216 2851 2228
rect 2849 2204 2853 2216
rect 2871 2204 2875 2236
rect 2881 2204 2885 2262
rect 2901 2224 2905 2261
rect 2965 2224 2969 2301
rect 2992 2259 2996 2316
rect 3000 2312 3004 2316
rect 3070 2313 3074 2356
rect 3000 2304 3018 2312
rect 3014 2293 3018 2304
rect 3067 2301 3074 2313
rect 2985 2247 2994 2259
rect 2985 2224 2989 2247
rect 3014 2236 3018 2281
rect 3005 2229 3018 2236
rect 3005 2224 3009 2229
rect 3065 2224 3069 2301
rect 3092 2259 3096 2316
rect 3100 2312 3104 2316
rect 3156 2312 3160 2316
rect 3100 2304 3118 2312
rect 3114 2293 3118 2304
rect 3142 2304 3160 2312
rect 3142 2293 3146 2304
rect 3085 2247 3094 2259
rect 3085 2224 3089 2247
rect 3114 2236 3118 2281
rect 3105 2229 3118 2236
rect 3142 2236 3146 2281
rect 3164 2259 3168 2316
rect 3186 2313 3190 2356
rect 3273 2353 3277 2376
rect 3269 2346 3277 2353
rect 3269 2317 3273 2346
rect 3281 2336 3285 2376
rect 3301 2324 3305 2356
rect 3309 2352 3313 2356
rect 3309 2350 3345 2352
rect 3309 2348 3333 2350
rect 3186 2301 3193 2313
rect 3251 2304 3255 2316
rect 3269 2311 3277 2317
rect 3166 2247 3175 2259
rect 3142 2229 3155 2236
rect 3105 2224 3109 2229
rect 3151 2224 3155 2229
rect 3171 2224 3175 2247
rect 3191 2224 3195 2301
rect 3251 2292 3253 2304
rect 3251 2224 3255 2292
rect 3273 2265 3277 2311
rect 3273 2204 3277 2253
rect 3301 2229 3307 2324
rect 3283 2225 3307 2229
rect 3283 2204 3287 2225
rect 3303 2220 3321 2221
rect 3303 2216 3333 2220
rect 3303 2204 3307 2216
rect 3341 2212 3345 2338
rect 3355 2330 3359 2356
rect 3375 2350 3379 2356
rect 3311 2208 3345 2212
rect 3311 2204 3315 2208
rect 3357 2204 3361 2318
rect 3373 2228 3377 2338
rect 3387 2316 3391 2356
rect 3382 2304 3385 2316
rect 3382 2240 3386 2304
rect 3407 2297 3411 2356
rect 3402 2289 3411 2297
rect 3402 2260 3406 2289
rect 3421 2274 3425 2356
rect 3441 2273 3445 2316
rect 3510 2313 3514 2356
rect 3507 2301 3514 2313
rect 3382 2236 3415 2240
rect 3381 2216 3383 2228
rect 3379 2204 3383 2216
rect 3389 2216 3391 2228
rect 3389 2204 3393 2216
rect 3411 2204 3415 2236
rect 3421 2204 3425 2262
rect 3441 2224 3445 2261
rect 3505 2224 3509 2301
rect 3532 2259 3536 2316
rect 3540 2312 3544 2316
rect 3540 2304 3558 2312
rect 3554 2293 3558 2304
rect 3617 2293 3621 2316
rect 3606 2281 3621 2293
rect 3625 2293 3629 2316
rect 3671 2312 3675 2316
rect 3662 2307 3675 2312
rect 3625 2281 3634 2293
rect 3525 2247 3534 2259
rect 3525 2224 3529 2247
rect 3554 2236 3558 2281
rect 3545 2229 3558 2236
rect 3545 2224 3549 2229
rect 3605 2204 3609 2281
rect 3625 2204 3629 2281
rect 3662 2273 3666 2307
rect 3681 2293 3685 2316
rect 3701 2311 3705 2316
rect 3662 2216 3666 2261
rect 3681 2217 3685 2281
rect 3785 2279 3789 2356
rect 3786 2267 3789 2279
rect 3783 2251 3789 2267
rect 3805 2279 3809 2356
rect 3865 2293 3869 2316
rect 3866 2281 3869 2293
rect 3805 2267 3814 2279
rect 3805 2251 3811 2267
rect 3783 2244 3797 2251
rect 3705 2232 3715 2244
rect 3711 2224 3715 2232
rect 3793 2224 3797 2244
rect 3803 2244 3811 2251
rect 3803 2224 3807 2244
rect 3860 2233 3866 2281
rect 3885 2259 3889 2316
rect 3905 2294 3909 2316
rect 3925 2294 3929 2316
rect 3905 2288 3918 2294
rect 3925 2293 3945 2294
rect 3985 2293 3989 2316
rect 3925 2288 3933 2293
rect 3914 2259 3918 2288
rect 3986 2281 3989 2293
rect 3887 2247 3889 2259
rect 3885 2245 3889 2247
rect 3885 2238 3898 2245
rect 3860 2229 3890 2233
rect 3886 2224 3890 2229
rect 3894 2224 3898 2238
rect 3914 2224 3918 2247
rect 3933 2239 3939 2281
rect 3922 2232 3939 2239
rect 3980 2233 3986 2281
rect 4005 2259 4009 2316
rect 4025 2294 4029 2316
rect 4045 2294 4049 2316
rect 4025 2288 4038 2294
rect 4045 2293 4065 2294
rect 4045 2288 4053 2293
rect 4034 2259 4038 2288
rect 4007 2247 4009 2259
rect 4005 2245 4009 2247
rect 4005 2238 4018 2245
rect 3922 2224 3926 2232
rect 3980 2229 4010 2233
rect 4006 2224 4010 2229
rect 4014 2224 4018 2238
rect 4034 2224 4038 2247
rect 4053 2239 4059 2281
rect 4095 2273 4099 2316
rect 4115 2274 4119 2356
rect 4129 2297 4133 2356
rect 4149 2316 4153 2356
rect 4161 2350 4165 2356
rect 4155 2304 4158 2316
rect 4129 2289 4138 2297
rect 4042 2232 4059 2239
rect 4042 2224 4046 2232
rect 4095 2224 4099 2261
rect 3662 2211 3675 2216
rect 3681 2211 3695 2217
rect 3671 2204 3675 2211
rect 3691 2204 3695 2211
rect 4115 2204 4119 2262
rect 4134 2260 4138 2289
rect 4154 2240 4158 2304
rect 4125 2236 4158 2240
rect 4125 2204 4129 2236
rect 4163 2228 4167 2338
rect 4181 2330 4185 2356
rect 4227 2352 4231 2356
rect 4195 2350 4231 2352
rect 4207 2348 4231 2350
rect 4149 2216 4151 2228
rect 4147 2204 4151 2216
rect 4157 2216 4159 2228
rect 4157 2204 4161 2216
rect 4179 2204 4183 2318
rect 4195 2212 4199 2338
rect 4235 2324 4239 2356
rect 4255 2336 4259 2376
rect 4263 2353 4267 2376
rect 4263 2346 4271 2353
rect 4233 2229 4239 2324
rect 4267 2317 4271 2346
rect 4263 2311 4271 2317
rect 4353 2353 4357 2376
rect 4349 2346 4357 2353
rect 4349 2317 4353 2346
rect 4361 2336 4365 2376
rect 4381 2324 4385 2356
rect 4389 2352 4393 2356
rect 4389 2350 4425 2352
rect 4389 2348 4413 2350
rect 4263 2265 4267 2311
rect 4285 2304 4289 2316
rect 4287 2292 4289 2304
rect 4233 2225 4257 2229
rect 4219 2220 4237 2221
rect 4207 2216 4237 2220
rect 4195 2208 4229 2212
rect 4225 2204 4229 2208
rect 4233 2204 4237 2216
rect 4253 2204 4257 2225
rect 4263 2204 4267 2253
rect 4285 2224 4289 2292
rect 4331 2304 4335 2316
rect 4349 2311 4357 2317
rect 4331 2292 4333 2304
rect 4331 2224 4335 2292
rect 4353 2265 4357 2311
rect 4353 2204 4357 2253
rect 4381 2229 4387 2324
rect 4363 2225 4387 2229
rect 4363 2204 4367 2225
rect 4383 2220 4401 2221
rect 4383 2216 4413 2220
rect 4383 2204 4387 2216
rect 4421 2212 4425 2338
rect 4435 2330 4439 2356
rect 4455 2350 4459 2356
rect 4391 2208 4425 2212
rect 4391 2204 4395 2208
rect 4437 2204 4441 2318
rect 4453 2228 4457 2338
rect 4467 2316 4471 2356
rect 4462 2304 4465 2316
rect 4462 2240 4466 2304
rect 4487 2297 4491 2356
rect 4482 2289 4491 2297
rect 4482 2260 4486 2289
rect 4501 2274 4505 2356
rect 4521 2273 4525 2316
rect 4576 2312 4580 2316
rect 4562 2304 4580 2312
rect 4562 2293 4566 2304
rect 4462 2236 4495 2240
rect 4461 2216 4463 2228
rect 4459 2204 4463 2216
rect 4469 2216 4471 2228
rect 4469 2204 4473 2216
rect 4491 2204 4495 2236
rect 4501 2204 4505 2262
rect 4521 2224 4525 2261
rect 4562 2236 4566 2281
rect 4584 2259 4588 2316
rect 4606 2313 4610 2356
rect 4606 2301 4613 2313
rect 4586 2247 4595 2259
rect 4562 2229 4575 2236
rect 4571 2224 4575 2229
rect 4591 2224 4595 2247
rect 4611 2224 4615 2301
rect 4671 2279 4675 2356
rect 4666 2267 4675 2279
rect 4669 2251 4675 2267
rect 4691 2279 4695 2356
rect 4691 2267 4694 2279
rect 4691 2251 4697 2267
rect 4669 2244 4677 2251
rect 4673 2224 4677 2244
rect 4683 2244 4697 2251
rect 4683 2224 4687 2244
rect 68 2180 72 2184
rect 76 2180 80 2184
rect 84 2180 88 2184
rect 145 2180 149 2184
rect 165 2180 169 2184
rect 185 2180 189 2184
rect 231 2180 235 2184
rect 251 2180 255 2184
rect 271 2180 275 2184
rect 332 2180 336 2184
rect 340 2180 344 2184
rect 348 2180 352 2184
rect 434 2180 438 2184
rect 442 2180 446 2184
rect 464 2180 468 2184
rect 531 2180 535 2184
rect 551 2180 555 2184
rect 571 2180 575 2184
rect 652 2180 656 2184
rect 674 2180 678 2184
rect 682 2180 686 2184
rect 731 2180 735 2184
rect 815 2180 819 2184
rect 835 2180 839 2184
rect 845 2180 849 2184
rect 893 2180 897 2184
rect 903 2180 907 2184
rect 971 2180 975 2184
rect 981 2180 985 2184
rect 1001 2180 1005 2184
rect 1085 2180 1089 2184
rect 1105 2180 1109 2184
rect 1125 2180 1129 2184
rect 1185 2180 1189 2184
rect 1205 2180 1209 2184
rect 1225 2180 1229 2184
rect 1275 2180 1279 2184
rect 1295 2180 1299 2184
rect 1305 2180 1309 2184
rect 1327 2180 1331 2184
rect 1337 2180 1341 2184
rect 1359 2180 1363 2184
rect 1405 2180 1409 2184
rect 1413 2180 1417 2184
rect 1433 2180 1437 2184
rect 1443 2180 1447 2184
rect 1465 2180 1469 2184
rect 1525 2180 1529 2184
rect 1545 2180 1549 2184
rect 1565 2180 1569 2184
rect 1615 2180 1619 2184
rect 1635 2180 1639 2184
rect 1645 2180 1649 2184
rect 1667 2180 1671 2184
rect 1677 2180 1681 2184
rect 1699 2180 1703 2184
rect 1745 2180 1749 2184
rect 1753 2180 1757 2184
rect 1773 2180 1777 2184
rect 1783 2180 1787 2184
rect 1805 2180 1809 2184
rect 1865 2180 1869 2184
rect 1925 2180 1929 2184
rect 1971 2180 1975 2184
rect 1991 2180 1995 2184
rect 2011 2180 2015 2184
rect 2075 2180 2079 2184
rect 2095 2180 2099 2184
rect 2105 2180 2109 2184
rect 2127 2180 2131 2184
rect 2137 2180 2141 2184
rect 2159 2180 2163 2184
rect 2205 2180 2209 2184
rect 2213 2180 2217 2184
rect 2233 2180 2237 2184
rect 2243 2180 2247 2184
rect 2265 2180 2269 2184
rect 2332 2180 2336 2184
rect 2354 2180 2358 2184
rect 2362 2180 2366 2184
rect 2432 2180 2436 2184
rect 2454 2180 2458 2184
rect 2462 2180 2466 2184
rect 2512 2180 2516 2184
rect 2520 2180 2524 2184
rect 2528 2180 2532 2184
rect 2611 2180 2615 2184
rect 2621 2180 2625 2184
rect 2641 2180 2645 2184
rect 2711 2180 2715 2184
rect 2733 2180 2737 2184
rect 2743 2180 2747 2184
rect 2763 2180 2767 2184
rect 2771 2180 2775 2184
rect 2817 2180 2821 2184
rect 2839 2180 2843 2184
rect 2849 2180 2853 2184
rect 2871 2180 2875 2184
rect 2881 2180 2885 2184
rect 2901 2180 2905 2184
rect 2965 2180 2969 2184
rect 2985 2180 2989 2184
rect 3005 2180 3009 2184
rect 3065 2180 3069 2184
rect 3085 2180 3089 2184
rect 3105 2180 3109 2184
rect 3151 2180 3155 2184
rect 3171 2180 3175 2184
rect 3191 2180 3195 2184
rect 3251 2180 3255 2184
rect 3273 2180 3277 2184
rect 3283 2180 3287 2184
rect 3303 2180 3307 2184
rect 3311 2180 3315 2184
rect 3357 2180 3361 2184
rect 3379 2180 3383 2184
rect 3389 2180 3393 2184
rect 3411 2180 3415 2184
rect 3421 2180 3425 2184
rect 3441 2180 3445 2184
rect 3505 2180 3509 2184
rect 3525 2180 3529 2184
rect 3545 2180 3549 2184
rect 3605 2180 3609 2184
rect 3625 2180 3629 2184
rect 3671 2180 3675 2184
rect 3691 2180 3695 2184
rect 3711 2180 3715 2184
rect 3793 2180 3797 2184
rect 3803 2180 3807 2184
rect 3886 2180 3890 2184
rect 3894 2180 3898 2184
rect 3914 2180 3918 2184
rect 3922 2180 3926 2184
rect 4006 2180 4010 2184
rect 4014 2180 4018 2184
rect 4034 2180 4038 2184
rect 4042 2180 4046 2184
rect 4095 2180 4099 2184
rect 4115 2180 4119 2184
rect 4125 2180 4129 2184
rect 4147 2180 4151 2184
rect 4157 2180 4161 2184
rect 4179 2180 4183 2184
rect 4225 2180 4229 2184
rect 4233 2180 4237 2184
rect 4253 2180 4257 2184
rect 4263 2180 4267 2184
rect 4285 2180 4289 2184
rect 4331 2180 4335 2184
rect 4353 2180 4357 2184
rect 4363 2180 4367 2184
rect 4383 2180 4387 2184
rect 4391 2180 4395 2184
rect 4437 2180 4441 2184
rect 4459 2180 4463 2184
rect 4469 2180 4473 2184
rect 4491 2180 4495 2184
rect 4501 2180 4505 2184
rect 4521 2180 4525 2184
rect 4571 2180 4575 2184
rect 4591 2180 4595 2184
rect 4611 2180 4615 2184
rect 4673 2180 4677 2184
rect 4683 2180 4687 2184
rect 43 2156 47 2160
rect 65 2156 69 2160
rect 125 2156 129 2160
rect 145 2156 149 2160
rect 165 2156 169 2160
rect 248 2156 252 2160
rect 256 2156 260 2160
rect 264 2156 268 2160
rect 314 2156 318 2160
rect 322 2156 326 2160
rect 344 2156 348 2160
rect 414 2156 418 2160
rect 422 2156 426 2160
rect 444 2156 448 2160
rect 512 2156 516 2160
rect 520 2156 524 2160
rect 528 2156 532 2160
rect 612 2156 616 2160
rect 620 2156 624 2160
rect 628 2156 632 2160
rect 714 2156 718 2160
rect 722 2156 726 2160
rect 744 2156 748 2160
rect 825 2156 829 2160
rect 845 2156 849 2160
rect 865 2156 869 2160
rect 912 2156 916 2160
rect 920 2156 924 2160
rect 928 2156 932 2160
rect 1012 2156 1016 2160
rect 1020 2156 1024 2160
rect 1028 2156 1032 2160
rect 1112 2156 1116 2160
rect 1120 2156 1124 2160
rect 1128 2156 1132 2160
rect 1214 2156 1218 2160
rect 1222 2156 1226 2160
rect 1244 2156 1248 2160
rect 1311 2156 1315 2160
rect 1331 2156 1335 2160
rect 1413 2156 1417 2160
rect 1423 2156 1427 2160
rect 1493 2156 1497 2160
rect 1503 2156 1507 2160
rect 1553 2156 1557 2160
rect 1563 2156 1567 2160
rect 1645 2156 1649 2160
rect 1665 2156 1669 2160
rect 1685 2156 1689 2160
rect 1734 2156 1738 2160
rect 1742 2156 1746 2160
rect 1764 2156 1768 2160
rect 1831 2156 1835 2160
rect 1851 2156 1855 2160
rect 1925 2156 1929 2160
rect 1945 2156 1949 2160
rect 1965 2156 1969 2160
rect 2011 2156 2015 2160
rect 2031 2156 2035 2160
rect 2051 2156 2055 2160
rect 2125 2156 2129 2160
rect 2145 2156 2149 2160
rect 2165 2156 2169 2160
rect 2225 2156 2229 2160
rect 2245 2156 2249 2160
rect 2265 2156 2269 2160
rect 2285 2156 2289 2160
rect 2305 2156 2309 2160
rect 2325 2156 2329 2160
rect 2345 2156 2349 2160
rect 2365 2156 2369 2160
rect 2413 2156 2417 2160
rect 2423 2156 2427 2160
rect 2515 2156 2519 2160
rect 2535 2156 2539 2160
rect 2545 2156 2549 2160
rect 2591 2156 2595 2160
rect 2611 2156 2615 2160
rect 2631 2156 2635 2160
rect 2713 2156 2717 2160
rect 2723 2156 2727 2160
rect 2773 2156 2777 2160
rect 2783 2156 2787 2160
rect 2855 2156 2859 2160
rect 2875 2156 2879 2160
rect 2885 2156 2889 2160
rect 2907 2156 2911 2160
rect 2917 2156 2921 2160
rect 2939 2156 2943 2160
rect 2985 2156 2989 2160
rect 2993 2156 2997 2160
rect 3013 2156 3017 2160
rect 3023 2156 3027 2160
rect 3045 2156 3049 2160
rect 3112 2156 3116 2160
rect 3134 2156 3138 2160
rect 3142 2156 3146 2160
rect 3191 2156 3195 2160
rect 3211 2156 3215 2160
rect 3306 2156 3310 2160
rect 3314 2156 3318 2160
rect 3334 2156 3338 2160
rect 3342 2156 3346 2160
rect 3395 2156 3399 2160
rect 3415 2156 3419 2160
rect 3425 2156 3429 2160
rect 3447 2156 3451 2160
rect 3457 2156 3461 2160
rect 3479 2156 3483 2160
rect 3525 2156 3529 2160
rect 3533 2156 3537 2160
rect 3553 2156 3557 2160
rect 3563 2156 3567 2160
rect 3585 2156 3589 2160
rect 3631 2156 3635 2160
rect 3651 2156 3655 2160
rect 3671 2156 3675 2160
rect 3735 2156 3739 2160
rect 3755 2156 3759 2160
rect 3765 2156 3769 2160
rect 3787 2156 3791 2160
rect 3797 2156 3801 2160
rect 3819 2156 3823 2160
rect 3865 2156 3869 2160
rect 3873 2156 3877 2160
rect 3893 2156 3897 2160
rect 3903 2156 3907 2160
rect 3925 2156 3929 2160
rect 3971 2156 3975 2160
rect 3993 2156 3997 2160
rect 4003 2156 4007 2160
rect 4023 2156 4027 2160
rect 4031 2156 4035 2160
rect 4077 2156 4081 2160
rect 4099 2156 4103 2160
rect 4109 2156 4113 2160
rect 4131 2156 4135 2160
rect 4141 2156 4145 2160
rect 4161 2156 4165 2160
rect 4246 2156 4250 2160
rect 4254 2156 4258 2160
rect 4274 2156 4278 2160
rect 4282 2156 4286 2160
rect 4331 2156 4335 2160
rect 4405 2156 4409 2160
rect 4425 2156 4429 2160
rect 4485 2156 4489 2160
rect 4505 2156 4509 2160
rect 4551 2156 4555 2160
rect 4573 2156 4577 2160
rect 4583 2156 4587 2160
rect 4603 2156 4607 2160
rect 4611 2156 4615 2160
rect 4657 2156 4661 2160
rect 4679 2156 4683 2160
rect 4689 2156 4693 2160
rect 4711 2156 4715 2160
rect 4721 2156 4725 2160
rect 4741 2156 4745 2160
rect 43 2110 47 2116
rect 43 2098 45 2110
rect 65 2059 69 2136
rect 65 2047 74 2059
rect 43 2030 45 2042
rect 43 2024 47 2030
rect 65 1984 69 2047
rect 125 2039 129 2116
rect 145 2093 149 2116
rect 165 2111 169 2116
rect 165 2104 178 2111
rect 145 2081 154 2093
rect 127 2027 134 2039
rect 130 1984 134 2027
rect 152 2024 156 2081
rect 174 2059 178 2104
rect 314 2112 318 2116
rect 299 2106 318 2112
rect 174 2036 178 2047
rect 248 2039 252 2096
rect 160 2028 178 2036
rect 160 2024 164 2028
rect 225 2027 233 2039
rect 245 2027 252 2039
rect 225 1984 229 2027
rect 256 2019 260 2096
rect 264 2039 268 2096
rect 299 2093 306 2106
rect 299 2044 306 2081
rect 322 2079 326 2116
rect 344 2093 348 2136
rect 414 2112 418 2116
rect 399 2106 418 2112
rect 399 2093 406 2106
rect 346 2081 355 2093
rect 320 2044 326 2067
rect 264 2027 274 2039
rect 299 2038 315 2044
rect 320 2038 335 2044
rect 254 2000 260 2007
rect 245 1996 260 2000
rect 274 1996 280 2027
rect 311 2024 315 2038
rect 331 2024 335 2038
rect 351 2024 355 2081
rect 399 2044 406 2081
rect 422 2079 426 2116
rect 444 2093 448 2136
rect 714 2112 718 2116
rect 699 2106 718 2112
rect 446 2081 455 2093
rect 420 2044 426 2067
rect 399 2038 415 2044
rect 420 2038 435 2044
rect 411 2024 415 2038
rect 431 2024 435 2038
rect 451 2024 455 2081
rect 512 2039 516 2096
rect 506 2027 516 2039
rect 245 1984 249 1996
rect 265 1992 280 1996
rect 265 1984 269 1992
rect 500 1996 506 2027
rect 520 2019 524 2096
rect 528 2039 532 2096
rect 612 2039 616 2096
rect 528 2027 535 2039
rect 547 2027 555 2039
rect 606 2027 616 2039
rect 520 2000 526 2007
rect 520 1996 535 2000
rect 500 1992 515 1996
rect 511 1984 515 1992
rect 531 1984 535 1996
rect 551 1984 555 2027
rect 600 1996 606 2027
rect 620 2019 624 2096
rect 628 2039 632 2096
rect 699 2093 706 2106
rect 699 2044 706 2081
rect 722 2079 726 2116
rect 744 2093 748 2136
rect 746 2081 755 2093
rect 720 2044 726 2067
rect 628 2027 635 2039
rect 647 2027 655 2039
rect 699 2038 715 2044
rect 720 2038 735 2044
rect 620 2000 626 2007
rect 620 1996 635 2000
rect 600 1992 615 1996
rect 611 1984 615 1992
rect 631 1984 635 1996
rect 651 1984 655 2027
rect 711 2024 715 2038
rect 731 2024 735 2038
rect 751 2024 755 2081
rect 825 2039 829 2116
rect 845 2093 849 2116
rect 865 2111 869 2116
rect 865 2104 878 2111
rect 845 2081 854 2093
rect 827 2027 834 2039
rect 830 1984 834 2027
rect 852 2024 856 2081
rect 874 2059 878 2104
rect 1214 2112 1218 2116
rect 1199 2106 1218 2112
rect 874 2036 878 2047
rect 912 2039 916 2096
rect 860 2028 878 2036
rect 860 2024 864 2028
rect 906 2027 916 2039
rect 900 1996 906 2027
rect 920 2019 924 2096
rect 928 2039 932 2096
rect 1012 2039 1016 2096
rect 928 2027 935 2039
rect 947 2027 955 2039
rect 1006 2027 1016 2039
rect 920 2000 926 2007
rect 920 1996 935 2000
rect 900 1992 915 1996
rect 911 1984 915 1992
rect 931 1984 935 1996
rect 951 1984 955 2027
rect 1000 1996 1006 2027
rect 1020 2019 1024 2096
rect 1028 2039 1032 2096
rect 1112 2039 1116 2096
rect 1028 2027 1035 2039
rect 1047 2027 1055 2039
rect 1106 2027 1116 2039
rect 1020 2000 1026 2007
rect 1020 1996 1035 2000
rect 1000 1992 1015 1996
rect 1011 1984 1015 1992
rect 1031 1984 1035 1996
rect 1051 1984 1055 2027
rect 1100 1996 1106 2027
rect 1120 2019 1124 2096
rect 1128 2039 1132 2096
rect 1199 2093 1206 2106
rect 1199 2044 1206 2081
rect 1222 2079 1226 2116
rect 1244 2093 1248 2136
rect 1246 2081 1255 2093
rect 1220 2044 1226 2067
rect 1128 2027 1135 2039
rect 1147 2027 1155 2039
rect 1199 2038 1215 2044
rect 1220 2038 1235 2044
rect 1120 2000 1126 2007
rect 1120 1996 1135 2000
rect 1100 1992 1115 1996
rect 1111 1984 1115 1992
rect 1131 1984 1135 1996
rect 1151 1984 1155 2027
rect 1211 2024 1215 2038
rect 1231 2024 1235 2038
rect 1251 2024 1255 2081
rect 1311 2059 1315 2136
rect 1331 2059 1335 2136
rect 1413 2096 1417 2116
rect 1403 2089 1417 2096
rect 1423 2096 1427 2116
rect 1493 2096 1497 2116
rect 1423 2089 1431 2096
rect 1403 2073 1409 2089
rect 1406 2061 1409 2073
rect 1306 2047 1315 2059
rect 1311 2024 1315 2047
rect 1319 2047 1334 2059
rect 1319 2024 1323 2047
rect 1405 1984 1409 2061
rect 1425 2073 1431 2089
rect 1483 2089 1497 2096
rect 1503 2096 1507 2116
rect 1553 2096 1557 2116
rect 1503 2089 1511 2096
rect 1483 2073 1489 2089
rect 1425 2061 1434 2073
rect 1486 2061 1489 2073
rect 1425 1984 1429 2061
rect 1485 1984 1489 2061
rect 1505 2073 1511 2089
rect 1549 2089 1557 2096
rect 1563 2096 1567 2116
rect 1563 2089 1577 2096
rect 1549 2073 1555 2089
rect 1505 2061 1514 2073
rect 1546 2061 1555 2073
rect 1505 1984 1509 2061
rect 1551 1984 1555 2061
rect 1571 2073 1577 2089
rect 1571 2061 1574 2073
rect 1571 1984 1575 2061
rect 1645 2039 1649 2116
rect 1665 2093 1669 2116
rect 1685 2111 1689 2116
rect 1734 2112 1738 2116
rect 1685 2104 1698 2111
rect 1665 2081 1674 2093
rect 1647 2027 1654 2039
rect 1650 1984 1654 2027
rect 1672 2024 1676 2081
rect 1694 2059 1698 2104
rect 1719 2106 1738 2112
rect 1719 2093 1726 2106
rect 1694 2036 1698 2047
rect 1719 2044 1726 2081
rect 1742 2079 1746 2116
rect 1764 2093 1768 2136
rect 1766 2081 1775 2093
rect 1740 2044 1746 2067
rect 1719 2038 1735 2044
rect 1740 2038 1755 2044
rect 1680 2028 1698 2036
rect 1680 2024 1684 2028
rect 1731 2024 1735 2038
rect 1751 2024 1755 2038
rect 1771 2024 1775 2081
rect 1831 2059 1835 2136
rect 1851 2059 1855 2136
rect 2591 2129 2595 2136
rect 2611 2129 2615 2136
rect 2582 2124 2595 2129
rect 1826 2047 1835 2059
rect 1831 2024 1835 2047
rect 1839 2047 1854 2059
rect 1839 2024 1843 2047
rect 1925 2039 1929 2116
rect 1945 2093 1949 2116
rect 1965 2111 1969 2116
rect 2011 2111 2015 2116
rect 1965 2104 1978 2111
rect 1945 2081 1954 2093
rect 1927 2027 1934 2039
rect 1930 1984 1934 2027
rect 1952 2024 1956 2081
rect 1974 2059 1978 2104
rect 2002 2104 2015 2111
rect 2002 2059 2006 2104
rect 2031 2093 2035 2116
rect 2026 2081 2035 2093
rect 1974 2036 1978 2047
rect 1960 2028 1978 2036
rect 2002 2036 2006 2047
rect 2002 2028 2020 2036
rect 1960 2024 1964 2028
rect 2016 2024 2020 2028
rect 2024 2024 2028 2081
rect 2051 2039 2055 2116
rect 2125 2039 2129 2116
rect 2145 2093 2149 2116
rect 2165 2111 2169 2116
rect 2165 2104 2178 2111
rect 2145 2081 2154 2093
rect 2046 2027 2053 2039
rect 2127 2027 2134 2039
rect 2046 1984 2050 2027
rect 2130 1984 2134 2027
rect 2152 2024 2156 2081
rect 2174 2059 2178 2104
rect 2225 2096 2229 2116
rect 2245 2096 2249 2116
rect 2265 2096 2269 2116
rect 2285 2096 2289 2116
rect 2305 2096 2309 2116
rect 2325 2096 2329 2116
rect 2225 2084 2238 2096
rect 2265 2084 2278 2096
rect 2305 2084 2318 2096
rect 2345 2093 2349 2116
rect 2365 2093 2369 2116
rect 2413 2096 2417 2116
rect 2174 2036 2178 2047
rect 2160 2028 2178 2036
rect 2160 2024 2164 2028
rect 2225 2024 2229 2084
rect 2245 2024 2249 2084
rect 2265 2024 2269 2084
rect 2285 2024 2289 2084
rect 2305 2024 2309 2084
rect 2325 2024 2329 2084
rect 2345 2081 2354 2093
rect 2366 2081 2369 2093
rect 2345 2024 2349 2081
rect 2365 2024 2369 2081
rect 2409 2089 2417 2096
rect 2423 2096 2427 2116
rect 2515 2110 2519 2116
rect 2501 2098 2513 2110
rect 2423 2089 2437 2096
rect 2409 2073 2415 2089
rect 2406 2061 2415 2073
rect 2411 1984 2415 2061
rect 2431 2073 2437 2089
rect 2431 2061 2434 2073
rect 2431 1984 2435 2061
rect 2501 2024 2505 2098
rect 2535 2073 2539 2116
rect 2526 2061 2539 2073
rect 2523 1984 2527 2061
rect 2545 2059 2549 2116
rect 2582 2079 2586 2124
rect 2545 2047 2554 2059
rect 2545 1984 2549 2047
rect 2582 2033 2586 2067
rect 2601 2123 2615 2129
rect 2601 2059 2605 2123
rect 2631 2108 2635 2116
rect 2625 2096 2635 2108
rect 2713 2096 2717 2116
rect 2703 2089 2717 2096
rect 2723 2096 2727 2116
rect 2773 2096 2777 2116
rect 2723 2089 2731 2096
rect 2703 2073 2709 2089
rect 2706 2061 2709 2073
rect 2582 2028 2595 2033
rect 2591 2024 2595 2028
rect 2601 2024 2605 2047
rect 2621 2024 2625 2029
rect 2705 1984 2709 2061
rect 2725 2073 2731 2089
rect 2769 2089 2777 2096
rect 2783 2096 2787 2116
rect 2783 2089 2797 2096
rect 2769 2073 2775 2089
rect 2725 2061 2734 2073
rect 2766 2061 2775 2073
rect 2725 1984 2729 2061
rect 2771 1984 2775 2061
rect 2791 2073 2797 2089
rect 2855 2079 2859 2116
rect 2791 2061 2794 2073
rect 2875 2078 2879 2136
rect 2885 2104 2889 2136
rect 2907 2124 2911 2136
rect 2909 2112 2911 2124
rect 2917 2124 2921 2136
rect 2917 2112 2919 2124
rect 2885 2100 2918 2104
rect 2791 1984 2795 2061
rect 2855 2024 2859 2067
rect 2875 1984 2879 2066
rect 2894 2051 2898 2080
rect 2889 2043 2898 2051
rect 2889 1984 2893 2043
rect 2914 2036 2918 2100
rect 2915 2024 2918 2036
rect 2909 1984 2913 2024
rect 2923 2002 2927 2112
rect 2939 2022 2943 2136
rect 2985 2132 2989 2136
rect 2955 2128 2989 2132
rect 2921 1984 2925 1990
rect 2941 1984 2945 2010
rect 2955 2002 2959 2128
rect 2993 2124 2997 2136
rect 2967 2120 2997 2124
rect 2979 2119 2997 2120
rect 3013 2115 3017 2136
rect 2993 2111 3017 2115
rect 2993 2016 2999 2111
rect 3023 2087 3027 2136
rect 3023 2029 3027 2075
rect 3045 2048 3049 2116
rect 3112 2093 3116 2136
rect 3047 2036 3049 2048
rect 3023 2023 3031 2029
rect 3045 2024 3049 2036
rect 3105 2081 3114 2093
rect 3105 2024 3109 2081
rect 3134 2079 3138 2116
rect 3142 2112 3146 2116
rect 3142 2106 3161 2112
rect 3154 2093 3161 2106
rect 3134 2044 3140 2067
rect 3154 2044 3161 2081
rect 3191 2059 3195 2136
rect 3211 2059 3215 2136
rect 3306 2111 3310 2116
rect 3280 2107 3310 2111
rect 3280 2059 3286 2107
rect 3314 2102 3318 2116
rect 3305 2095 3318 2102
rect 3305 2093 3309 2095
rect 3334 2093 3338 2116
rect 3342 2108 3346 2116
rect 3342 2101 3359 2108
rect 3307 2081 3309 2093
rect 3186 2047 3195 2059
rect 3125 2038 3140 2044
rect 3145 2038 3161 2044
rect 3125 2024 3129 2038
rect 3145 2024 3149 2038
rect 3191 2024 3195 2047
rect 3199 2047 3214 2059
rect 3286 2047 3289 2059
rect 3199 2024 3203 2047
rect 3285 2024 3289 2047
rect 3305 2024 3309 2081
rect 3334 2052 3338 2081
rect 3353 2059 3359 2101
rect 3395 2079 3399 2116
rect 3415 2078 3419 2136
rect 3425 2104 3429 2136
rect 3447 2124 3451 2136
rect 3449 2112 3451 2124
rect 3457 2124 3461 2136
rect 3457 2112 3459 2124
rect 3425 2100 3458 2104
rect 3325 2046 3338 2052
rect 3345 2047 3353 2052
rect 3345 2046 3365 2047
rect 3325 2024 3329 2046
rect 3345 2024 3349 2046
rect 3395 2024 3399 2067
rect 2967 1990 2991 1992
rect 2955 1988 2991 1990
rect 2987 1984 2991 1988
rect 2995 1984 2999 2016
rect 3015 1964 3019 2004
rect 3027 1994 3031 2023
rect 3023 1987 3031 1994
rect 3023 1964 3027 1987
rect 3415 1984 3419 2066
rect 3434 2051 3438 2080
rect 3429 2043 3438 2051
rect 3429 1984 3433 2043
rect 3454 2036 3458 2100
rect 3455 2024 3458 2036
rect 3449 1984 3453 2024
rect 3463 2002 3467 2112
rect 3479 2022 3483 2136
rect 3525 2132 3529 2136
rect 3495 2128 3529 2132
rect 3461 1984 3465 1990
rect 3481 1984 3485 2010
rect 3495 2002 3499 2128
rect 3533 2124 3537 2136
rect 3507 2120 3537 2124
rect 3519 2119 3537 2120
rect 3553 2115 3557 2136
rect 3533 2111 3557 2115
rect 3533 2016 3539 2111
rect 3563 2087 3567 2136
rect 3563 2029 3567 2075
rect 3585 2048 3589 2116
rect 3631 2111 3635 2116
rect 3622 2104 3635 2111
rect 3622 2059 3626 2104
rect 3651 2093 3655 2116
rect 3646 2081 3655 2093
rect 3587 2036 3589 2048
rect 3563 2023 3571 2029
rect 3585 2024 3589 2036
rect 3622 2036 3626 2047
rect 3622 2028 3640 2036
rect 3636 2024 3640 2028
rect 3644 2024 3648 2081
rect 3671 2039 3675 2116
rect 3735 2079 3739 2116
rect 3755 2078 3759 2136
rect 3765 2104 3769 2136
rect 3787 2124 3791 2136
rect 3789 2112 3791 2124
rect 3797 2124 3801 2136
rect 3797 2112 3799 2124
rect 3765 2100 3798 2104
rect 3666 2027 3673 2039
rect 3507 1990 3531 1992
rect 3495 1988 3531 1990
rect 3527 1984 3531 1988
rect 3535 1984 3539 2016
rect 3555 1964 3559 2004
rect 3567 1994 3571 2023
rect 3563 1987 3571 1994
rect 3563 1964 3567 1987
rect 3666 1984 3670 2027
rect 3735 2024 3739 2067
rect 3755 1984 3759 2066
rect 3774 2051 3778 2080
rect 3769 2043 3778 2051
rect 3769 1984 3773 2043
rect 3794 2036 3798 2100
rect 3795 2024 3798 2036
rect 3789 1984 3793 2024
rect 3803 2002 3807 2112
rect 3819 2022 3823 2136
rect 3865 2132 3869 2136
rect 3835 2128 3869 2132
rect 3801 1984 3805 1990
rect 3821 1984 3825 2010
rect 3835 2002 3839 2128
rect 3873 2124 3877 2136
rect 3847 2120 3877 2124
rect 3859 2119 3877 2120
rect 3893 2115 3897 2136
rect 3873 2111 3897 2115
rect 3873 2016 3879 2111
rect 3903 2087 3907 2136
rect 3903 2029 3907 2075
rect 3925 2048 3929 2116
rect 3927 2036 3929 2048
rect 3903 2023 3911 2029
rect 3925 2024 3929 2036
rect 3971 2048 3975 2116
rect 3993 2087 3997 2136
rect 4003 2115 4007 2136
rect 4023 2124 4027 2136
rect 4031 2132 4035 2136
rect 4031 2128 4065 2132
rect 4023 2120 4053 2124
rect 4023 2119 4041 2120
rect 4003 2111 4027 2115
rect 3971 2036 3973 2048
rect 3971 2024 3975 2036
rect 3993 2029 3997 2075
rect 3847 1990 3871 1992
rect 3835 1988 3871 1990
rect 3867 1984 3871 1988
rect 3875 1984 3879 2016
rect 3895 1964 3899 2004
rect 3907 1994 3911 2023
rect 3903 1987 3911 1994
rect 3903 1964 3907 1987
rect 3989 2023 3997 2029
rect 3989 1994 3993 2023
rect 4021 2016 4027 2111
rect 3989 1987 3997 1994
rect 3993 1964 3997 1987
rect 4001 1964 4005 2004
rect 4021 1984 4025 2016
rect 4061 2002 4065 2128
rect 4077 2022 4081 2136
rect 4099 2124 4103 2136
rect 4101 2112 4103 2124
rect 4109 2124 4113 2136
rect 4109 2112 4111 2124
rect 4029 1990 4053 1992
rect 4029 1988 4065 1990
rect 4029 1984 4033 1988
rect 4075 1984 4079 2010
rect 4093 2002 4097 2112
rect 4131 2104 4135 2136
rect 4102 2100 4135 2104
rect 4102 2036 4106 2100
rect 4122 2051 4126 2080
rect 4141 2078 4145 2136
rect 4161 2079 4165 2116
rect 4246 2111 4250 2116
rect 4220 2107 4250 2111
rect 4122 2043 4131 2051
rect 4102 2024 4105 2036
rect 4095 1984 4099 1990
rect 4107 1984 4111 2024
rect 4127 1984 4131 2043
rect 4141 1984 4145 2066
rect 4161 2024 4165 2067
rect 4220 2059 4226 2107
rect 4254 2102 4258 2116
rect 4245 2095 4258 2102
rect 4245 2093 4249 2095
rect 4274 2093 4278 2116
rect 4282 2108 4286 2116
rect 4282 2101 4299 2108
rect 4247 2081 4249 2093
rect 4226 2047 4229 2059
rect 4225 2024 4229 2047
rect 4245 2024 4249 2081
rect 4274 2052 4278 2081
rect 4293 2059 4299 2101
rect 4331 2079 4335 2136
rect 4326 2067 4335 2079
rect 4265 2046 4278 2052
rect 4285 2047 4293 2052
rect 4285 2046 4305 2047
rect 4265 2024 4269 2046
rect 4285 2024 4289 2046
rect 4331 1984 4335 2067
rect 4405 2059 4409 2136
rect 4425 2059 4429 2136
rect 4485 2059 4489 2136
rect 4505 2059 4509 2136
rect 4406 2047 4421 2059
rect 4417 2024 4421 2047
rect 4425 2047 4434 2059
rect 4486 2047 4501 2059
rect 4425 2024 4429 2047
rect 4497 2024 4501 2047
rect 4505 2047 4514 2059
rect 4551 2048 4555 2116
rect 4573 2087 4577 2136
rect 4583 2115 4587 2136
rect 4603 2124 4607 2136
rect 4611 2132 4615 2136
rect 4611 2128 4645 2132
rect 4603 2120 4633 2124
rect 4603 2119 4621 2120
rect 4583 2111 4607 2115
rect 4505 2024 4509 2047
rect 4551 2036 4553 2048
rect 4551 2024 4555 2036
rect 4573 2029 4577 2075
rect 4569 2023 4577 2029
rect 4569 1994 4573 2023
rect 4601 2016 4607 2111
rect 4569 1987 4577 1994
rect 4573 1964 4577 1987
rect 4581 1964 4585 2004
rect 4601 1984 4605 2016
rect 4641 2002 4645 2128
rect 4657 2022 4661 2136
rect 4679 2124 4683 2136
rect 4681 2112 4683 2124
rect 4689 2124 4693 2136
rect 4689 2112 4691 2124
rect 4609 1990 4633 1992
rect 4609 1988 4645 1990
rect 4609 1984 4613 1988
rect 4655 1984 4659 2010
rect 4673 2002 4677 2112
rect 4711 2104 4715 2136
rect 4682 2100 4715 2104
rect 4682 2036 4686 2100
rect 4702 2051 4706 2080
rect 4721 2078 4725 2136
rect 4741 2079 4745 2116
rect 4702 2043 4711 2051
rect 4682 2024 4685 2036
rect 4675 1984 4679 1990
rect 4687 1984 4691 2024
rect 4707 1984 4711 2043
rect 4721 1984 4725 2066
rect 4741 2024 4745 2067
rect 43 1940 47 1944
rect 65 1940 69 1944
rect 130 1940 134 1944
rect 152 1940 156 1944
rect 160 1940 164 1944
rect 225 1940 229 1944
rect 245 1940 249 1944
rect 265 1940 269 1944
rect 311 1940 315 1944
rect 331 1940 335 1944
rect 351 1940 355 1944
rect 411 1940 415 1944
rect 431 1940 435 1944
rect 451 1940 455 1944
rect 511 1940 515 1944
rect 531 1940 535 1944
rect 551 1940 555 1944
rect 611 1940 615 1944
rect 631 1940 635 1944
rect 651 1940 655 1944
rect 711 1940 715 1944
rect 731 1940 735 1944
rect 751 1940 755 1944
rect 830 1940 834 1944
rect 852 1940 856 1944
rect 860 1940 864 1944
rect 911 1940 915 1944
rect 931 1940 935 1944
rect 951 1940 955 1944
rect 1011 1940 1015 1944
rect 1031 1940 1035 1944
rect 1051 1940 1055 1944
rect 1111 1940 1115 1944
rect 1131 1940 1135 1944
rect 1151 1940 1155 1944
rect 1211 1940 1215 1944
rect 1231 1940 1235 1944
rect 1251 1940 1255 1944
rect 1311 1940 1315 1944
rect 1319 1940 1323 1944
rect 1405 1940 1409 1944
rect 1425 1940 1429 1944
rect 1485 1940 1489 1944
rect 1505 1940 1509 1944
rect 1551 1940 1555 1944
rect 1571 1940 1575 1944
rect 1650 1940 1654 1944
rect 1672 1940 1676 1944
rect 1680 1940 1684 1944
rect 1731 1940 1735 1944
rect 1751 1940 1755 1944
rect 1771 1940 1775 1944
rect 1831 1940 1835 1944
rect 1839 1940 1843 1944
rect 1930 1940 1934 1944
rect 1952 1940 1956 1944
rect 1960 1940 1964 1944
rect 2016 1940 2020 1944
rect 2024 1940 2028 1944
rect 2046 1940 2050 1944
rect 2130 1940 2134 1944
rect 2152 1940 2156 1944
rect 2160 1940 2164 1944
rect 2225 1940 2229 1944
rect 2245 1940 2249 1944
rect 2265 1940 2269 1944
rect 2285 1940 2289 1944
rect 2305 1940 2309 1944
rect 2325 1940 2329 1944
rect 2345 1940 2349 1944
rect 2365 1940 2369 1944
rect 2411 1940 2415 1944
rect 2431 1940 2435 1944
rect 2501 1940 2505 1944
rect 2523 1940 2527 1944
rect 2545 1940 2549 1944
rect 2591 1940 2595 1944
rect 2601 1940 2605 1944
rect 2621 1940 2625 1944
rect 2705 1940 2709 1944
rect 2725 1940 2729 1944
rect 2771 1940 2775 1944
rect 2791 1940 2795 1944
rect 2855 1940 2859 1944
rect 2875 1940 2879 1944
rect 2889 1940 2893 1944
rect 2909 1940 2913 1944
rect 2921 1940 2925 1944
rect 2941 1940 2945 1944
rect 2987 1940 2991 1944
rect 2995 1940 2999 1944
rect 3015 1940 3019 1944
rect 3023 1940 3027 1944
rect 3045 1940 3049 1944
rect 3105 1940 3109 1944
rect 3125 1940 3129 1944
rect 3145 1940 3149 1944
rect 3191 1940 3195 1944
rect 3199 1940 3203 1944
rect 3285 1940 3289 1944
rect 3305 1940 3309 1944
rect 3325 1940 3329 1944
rect 3345 1940 3349 1944
rect 3395 1940 3399 1944
rect 3415 1940 3419 1944
rect 3429 1940 3433 1944
rect 3449 1940 3453 1944
rect 3461 1940 3465 1944
rect 3481 1940 3485 1944
rect 3527 1940 3531 1944
rect 3535 1940 3539 1944
rect 3555 1940 3559 1944
rect 3563 1940 3567 1944
rect 3585 1940 3589 1944
rect 3636 1940 3640 1944
rect 3644 1940 3648 1944
rect 3666 1940 3670 1944
rect 3735 1940 3739 1944
rect 3755 1940 3759 1944
rect 3769 1940 3773 1944
rect 3789 1940 3793 1944
rect 3801 1940 3805 1944
rect 3821 1940 3825 1944
rect 3867 1940 3871 1944
rect 3875 1940 3879 1944
rect 3895 1940 3899 1944
rect 3903 1940 3907 1944
rect 3925 1940 3929 1944
rect 3971 1940 3975 1944
rect 3993 1940 3997 1944
rect 4001 1940 4005 1944
rect 4021 1940 4025 1944
rect 4029 1940 4033 1944
rect 4075 1940 4079 1944
rect 4095 1940 4099 1944
rect 4107 1940 4111 1944
rect 4127 1940 4131 1944
rect 4141 1940 4145 1944
rect 4161 1940 4165 1944
rect 4225 1940 4229 1944
rect 4245 1940 4249 1944
rect 4265 1940 4269 1944
rect 4285 1940 4289 1944
rect 4331 1940 4335 1944
rect 4417 1940 4421 1944
rect 4425 1940 4429 1944
rect 4497 1940 4501 1944
rect 4505 1940 4509 1944
rect 4551 1940 4555 1944
rect 4573 1940 4577 1944
rect 4581 1940 4585 1944
rect 4601 1940 4605 1944
rect 4609 1940 4613 1944
rect 4655 1940 4659 1944
rect 4675 1940 4679 1944
rect 4687 1940 4691 1944
rect 4707 1940 4711 1944
rect 4721 1940 4725 1944
rect 4741 1940 4745 1944
rect 45 1916 49 1920
rect 65 1916 69 1920
rect 85 1916 89 1920
rect 105 1916 109 1920
rect 156 1916 160 1920
rect 164 1916 168 1920
rect 186 1916 190 1920
rect 251 1916 255 1920
rect 271 1916 275 1920
rect 345 1916 349 1920
rect 365 1916 369 1920
rect 385 1916 389 1920
rect 431 1916 435 1920
rect 451 1916 455 1920
rect 471 1916 475 1920
rect 491 1916 495 1920
rect 551 1916 555 1920
rect 573 1916 577 1920
rect 595 1916 599 1920
rect 665 1916 669 1920
rect 711 1916 715 1920
rect 733 1916 737 1920
rect 810 1916 814 1920
rect 832 1916 836 1920
rect 840 1916 844 1920
rect 896 1916 900 1920
rect 904 1916 908 1920
rect 926 1916 930 1920
rect 991 1916 995 1920
rect 1011 1916 1015 1920
rect 1031 1916 1035 1920
rect 1091 1916 1095 1920
rect 1151 1916 1155 1920
rect 1171 1916 1175 1920
rect 1191 1916 1195 1920
rect 1251 1916 1255 1920
rect 1271 1916 1275 1920
rect 1291 1916 1295 1920
rect 1365 1916 1369 1920
rect 1425 1916 1429 1920
rect 1445 1916 1449 1920
rect 1465 1916 1469 1920
rect 1485 1916 1489 1920
rect 1531 1916 1535 1920
rect 1551 1916 1555 1920
rect 1571 1916 1575 1920
rect 1631 1916 1635 1920
rect 1705 1916 1709 1920
rect 1765 1916 1769 1920
rect 1785 1916 1789 1920
rect 1805 1916 1809 1920
rect 1851 1916 1855 1920
rect 1873 1916 1877 1920
rect 1895 1916 1899 1920
rect 1955 1916 1959 1920
rect 1975 1916 1979 1920
rect 1989 1916 1993 1920
rect 2009 1916 2013 1920
rect 2021 1916 2025 1920
rect 2041 1916 2045 1920
rect 2087 1916 2091 1920
rect 2095 1916 2099 1920
rect 2115 1916 2119 1920
rect 2123 1916 2127 1920
rect 2145 1916 2149 1920
rect 2217 1916 2221 1920
rect 2225 1916 2229 1920
rect 2271 1916 2275 1920
rect 2336 1916 2340 1920
rect 2344 1916 2348 1920
rect 2366 1916 2370 1920
rect 2431 1916 2435 1920
rect 2439 1916 2443 1920
rect 2511 1916 2515 1920
rect 2519 1916 2523 1920
rect 2596 1916 2600 1920
rect 2604 1916 2608 1920
rect 2626 1916 2630 1920
rect 2705 1916 2709 1920
rect 2725 1916 2729 1920
rect 2797 1916 2801 1920
rect 2805 1916 2809 1920
rect 2856 1916 2860 1920
rect 2864 1916 2868 1920
rect 2886 1916 2890 1920
rect 2951 1916 2955 1920
rect 3037 1916 3041 1920
rect 3045 1916 3049 1920
rect 3091 1916 3095 1920
rect 3113 1916 3117 1920
rect 3121 1916 3125 1920
rect 3141 1916 3145 1920
rect 3149 1916 3153 1920
rect 3195 1916 3199 1920
rect 3215 1916 3219 1920
rect 3227 1916 3231 1920
rect 3247 1916 3251 1920
rect 3261 1916 3265 1920
rect 3281 1916 3285 1920
rect 3336 1916 3340 1920
rect 3344 1916 3348 1920
rect 3366 1916 3370 1920
rect 3431 1916 3435 1920
rect 3451 1916 3455 1920
rect 3511 1916 3515 1920
rect 3533 1916 3537 1920
rect 3541 1916 3545 1920
rect 3561 1916 3565 1920
rect 3569 1916 3573 1920
rect 3615 1916 3619 1920
rect 3635 1916 3639 1920
rect 3647 1916 3651 1920
rect 3667 1916 3671 1920
rect 3681 1916 3685 1920
rect 3701 1916 3705 1920
rect 3751 1916 3755 1920
rect 3773 1916 3777 1920
rect 3845 1916 3849 1920
rect 3865 1916 3869 1920
rect 3930 1916 3934 1920
rect 3952 1916 3956 1920
rect 3960 1916 3964 1920
rect 4030 1916 4034 1920
rect 4052 1916 4056 1920
rect 4060 1916 4064 1920
rect 4111 1916 4115 1920
rect 4121 1916 4125 1920
rect 4141 1916 4145 1920
rect 4225 1916 4229 1920
rect 4271 1916 4275 1920
rect 4291 1916 4295 1920
rect 4311 1916 4315 1920
rect 4397 1916 4401 1920
rect 4405 1916 4409 1920
rect 4451 1916 4455 1920
rect 4473 1916 4477 1920
rect 4481 1916 4485 1920
rect 4501 1916 4505 1920
rect 4509 1916 4513 1920
rect 4555 1916 4559 1920
rect 4575 1916 4579 1920
rect 4587 1916 4591 1920
rect 4607 1916 4611 1920
rect 4621 1916 4625 1920
rect 4641 1916 4645 1920
rect 4705 1916 4709 1920
rect 4725 1916 4729 1920
rect 45 1813 49 1836
rect 46 1801 49 1813
rect 40 1753 46 1801
rect 65 1779 69 1836
rect 85 1814 89 1836
rect 105 1814 109 1836
rect 156 1832 160 1836
rect 142 1824 160 1832
rect 85 1808 98 1814
rect 105 1813 125 1814
rect 142 1813 146 1824
rect 105 1808 113 1813
rect 94 1779 98 1808
rect 67 1767 69 1779
rect 65 1765 69 1767
rect 65 1758 78 1765
rect 40 1749 70 1753
rect 66 1744 70 1749
rect 74 1744 78 1758
rect 94 1744 98 1767
rect 113 1759 119 1801
rect 102 1752 119 1759
rect 142 1756 146 1801
rect 164 1779 168 1836
rect 186 1833 190 1876
rect 186 1821 193 1833
rect 166 1767 175 1779
rect 102 1744 106 1752
rect 142 1749 155 1756
rect 151 1744 155 1749
rect 171 1744 175 1767
rect 191 1744 195 1821
rect 251 1799 255 1876
rect 246 1787 255 1799
rect 249 1771 255 1787
rect 271 1799 275 1876
rect 345 1833 349 1876
rect 365 1864 369 1876
rect 385 1868 389 1876
rect 385 1864 400 1868
rect 365 1860 380 1864
rect 374 1853 380 1860
rect 345 1821 353 1833
rect 365 1821 372 1833
rect 271 1787 274 1799
rect 271 1771 277 1787
rect 249 1764 257 1771
rect 253 1744 257 1764
rect 263 1764 277 1771
rect 368 1764 372 1821
rect 376 1764 380 1841
rect 394 1833 400 1864
rect 384 1821 394 1833
rect 384 1764 388 1821
rect 431 1814 435 1836
rect 451 1814 455 1836
rect 415 1813 435 1814
rect 427 1808 435 1813
rect 442 1808 455 1814
rect 263 1744 267 1764
rect 421 1759 427 1801
rect 442 1779 446 1808
rect 471 1779 475 1836
rect 491 1813 495 1836
rect 551 1813 555 1876
rect 491 1801 494 1813
rect 546 1801 555 1813
rect 471 1767 473 1779
rect 421 1752 438 1759
rect 434 1744 438 1752
rect 442 1744 446 1767
rect 471 1765 475 1767
rect 462 1758 475 1765
rect 462 1744 466 1758
rect 494 1753 500 1801
rect 470 1749 500 1753
rect 470 1744 474 1749
rect 551 1744 555 1801
rect 573 1799 577 1876
rect 561 1787 574 1799
rect 561 1744 565 1787
rect 595 1762 599 1836
rect 587 1750 599 1762
rect 665 1779 669 1836
rect 711 1813 715 1876
rect 733 1830 737 1836
rect 810 1833 814 1876
rect 735 1818 737 1830
rect 807 1821 814 1833
rect 706 1801 715 1813
rect 665 1767 674 1779
rect 581 1744 585 1750
rect 665 1744 669 1767
rect 711 1724 715 1801
rect 735 1750 737 1762
rect 733 1744 737 1750
rect 805 1744 809 1821
rect 832 1779 836 1836
rect 840 1832 844 1836
rect 896 1832 900 1836
rect 840 1824 858 1832
rect 854 1813 858 1824
rect 882 1824 900 1832
rect 882 1813 886 1824
rect 825 1767 834 1779
rect 825 1744 829 1767
rect 854 1756 858 1801
rect 845 1749 858 1756
rect 882 1756 886 1801
rect 904 1779 908 1836
rect 926 1833 930 1876
rect 991 1868 995 1876
rect 980 1864 995 1868
rect 1011 1864 1015 1876
rect 980 1833 986 1864
rect 1000 1860 1015 1864
rect 1000 1853 1006 1860
rect 926 1821 933 1833
rect 986 1821 996 1833
rect 906 1767 915 1779
rect 882 1749 895 1756
rect 845 1744 849 1749
rect 891 1744 895 1749
rect 911 1744 915 1767
rect 931 1744 935 1821
rect 992 1764 996 1821
rect 1000 1764 1004 1841
rect 1031 1833 1035 1876
rect 1008 1821 1015 1833
rect 1027 1821 1035 1833
rect 1008 1764 1012 1821
rect 1091 1793 1095 1876
rect 1151 1868 1155 1876
rect 1140 1864 1155 1868
rect 1171 1864 1175 1876
rect 1140 1833 1146 1864
rect 1160 1860 1175 1864
rect 1160 1853 1166 1860
rect 1146 1821 1156 1833
rect 1086 1781 1095 1793
rect 1091 1724 1095 1781
rect 1152 1764 1156 1821
rect 1160 1764 1164 1841
rect 1191 1833 1195 1876
rect 1251 1868 1255 1876
rect 1240 1864 1255 1868
rect 1271 1864 1275 1876
rect 1240 1833 1246 1864
rect 1260 1860 1275 1864
rect 1260 1853 1266 1860
rect 1168 1821 1175 1833
rect 1187 1821 1195 1833
rect 1246 1821 1256 1833
rect 1168 1764 1172 1821
rect 1252 1764 1256 1821
rect 1260 1764 1264 1841
rect 1291 1833 1295 1876
rect 1268 1821 1275 1833
rect 1287 1821 1295 1833
rect 1268 1764 1272 1821
rect 1365 1793 1369 1876
rect 1531 1868 1535 1876
rect 1520 1864 1535 1868
rect 1551 1864 1555 1876
rect 1425 1813 1429 1836
rect 1426 1801 1429 1813
rect 1365 1781 1374 1793
rect 1365 1724 1369 1781
rect 1420 1753 1426 1801
rect 1445 1779 1449 1836
rect 1465 1814 1469 1836
rect 1485 1814 1489 1836
rect 1520 1833 1526 1864
rect 1540 1860 1555 1864
rect 1540 1853 1546 1860
rect 1526 1821 1536 1833
rect 1465 1808 1478 1814
rect 1485 1813 1505 1814
rect 1485 1808 1493 1813
rect 1474 1779 1478 1808
rect 1447 1767 1449 1779
rect 1445 1765 1449 1767
rect 1445 1758 1458 1765
rect 1420 1749 1450 1753
rect 1446 1744 1450 1749
rect 1454 1744 1458 1758
rect 1474 1744 1478 1767
rect 1493 1759 1499 1801
rect 1532 1764 1536 1821
rect 1540 1764 1544 1841
rect 1571 1833 1575 1876
rect 1548 1821 1555 1833
rect 1567 1821 1575 1833
rect 1548 1764 1552 1821
rect 1631 1793 1635 1876
rect 1626 1781 1635 1793
rect 1482 1752 1499 1759
rect 1482 1744 1486 1752
rect 1631 1724 1635 1781
rect 1705 1779 1709 1836
rect 1765 1833 1769 1876
rect 1785 1864 1789 1876
rect 1805 1868 1809 1876
rect 1805 1864 1820 1868
rect 1785 1860 1800 1864
rect 1794 1853 1800 1860
rect 1765 1821 1773 1833
rect 1785 1821 1792 1833
rect 1705 1767 1714 1779
rect 1705 1744 1709 1767
rect 1788 1764 1792 1821
rect 1796 1764 1800 1841
rect 1814 1833 1820 1864
rect 1804 1821 1814 1833
rect 1804 1764 1808 1821
rect 1851 1813 1855 1876
rect 1846 1801 1855 1813
rect 1851 1744 1855 1801
rect 1873 1799 1877 1876
rect 1861 1787 1874 1799
rect 1861 1744 1865 1787
rect 1895 1762 1899 1836
rect 1955 1793 1959 1836
rect 1975 1794 1979 1876
rect 1989 1817 1993 1876
rect 2009 1836 2013 1876
rect 2021 1870 2025 1876
rect 2015 1824 2018 1836
rect 1989 1809 1998 1817
rect 1887 1750 1899 1762
rect 1881 1744 1885 1750
rect 1955 1744 1959 1781
rect 1975 1724 1979 1782
rect 1994 1780 1998 1809
rect 2014 1760 2018 1824
rect 1985 1756 2018 1760
rect 1985 1724 1989 1756
rect 2023 1748 2027 1858
rect 2041 1850 2045 1876
rect 2087 1872 2091 1876
rect 2055 1870 2091 1872
rect 2067 1868 2091 1870
rect 2009 1736 2011 1748
rect 2007 1724 2011 1736
rect 2017 1736 2019 1748
rect 2017 1724 2021 1736
rect 2039 1724 2043 1838
rect 2055 1732 2059 1858
rect 2095 1844 2099 1876
rect 2115 1856 2119 1896
rect 2123 1873 2127 1896
rect 2123 1866 2131 1873
rect 2093 1749 2099 1844
rect 2127 1837 2131 1866
rect 2123 1831 2131 1837
rect 2123 1785 2127 1831
rect 2145 1824 2149 1836
rect 2147 1812 2149 1824
rect 2217 1813 2221 1836
rect 2093 1745 2117 1749
rect 2079 1740 2097 1741
rect 2067 1736 2097 1740
rect 2055 1728 2089 1732
rect 2085 1724 2089 1728
rect 2093 1724 2097 1736
rect 2113 1724 2117 1745
rect 2123 1724 2127 1773
rect 2145 1744 2149 1812
rect 2206 1801 2221 1813
rect 2225 1813 2229 1836
rect 2225 1801 2234 1813
rect 2205 1724 2209 1801
rect 2225 1724 2229 1801
rect 2271 1793 2275 1876
rect 2336 1832 2340 1836
rect 2322 1824 2340 1832
rect 2322 1813 2326 1824
rect 2266 1781 2275 1793
rect 2271 1724 2275 1781
rect 2322 1756 2326 1801
rect 2344 1779 2348 1836
rect 2366 1833 2370 1876
rect 2366 1821 2373 1833
rect 2346 1767 2355 1779
rect 2322 1749 2335 1756
rect 2331 1744 2335 1749
rect 2351 1744 2355 1767
rect 2371 1744 2375 1821
rect 2431 1813 2435 1836
rect 2426 1801 2435 1813
rect 2439 1813 2443 1836
rect 2511 1813 2515 1836
rect 2439 1801 2454 1813
rect 2506 1801 2515 1813
rect 2519 1813 2523 1836
rect 2596 1832 2600 1836
rect 2582 1824 2600 1832
rect 2582 1813 2586 1824
rect 2519 1801 2534 1813
rect 2431 1724 2435 1801
rect 2451 1724 2455 1801
rect 2511 1724 2515 1801
rect 2531 1724 2535 1801
rect 2582 1756 2586 1801
rect 2604 1779 2608 1836
rect 2626 1833 2630 1876
rect 2626 1821 2633 1833
rect 2606 1767 2615 1779
rect 2582 1749 2595 1756
rect 2591 1744 2595 1749
rect 2611 1744 2615 1767
rect 2631 1744 2635 1821
rect 2705 1799 2709 1876
rect 2706 1787 2709 1799
rect 2703 1771 2709 1787
rect 2725 1799 2729 1876
rect 2797 1813 2801 1836
rect 2786 1801 2801 1813
rect 2805 1813 2809 1836
rect 2856 1832 2860 1836
rect 2842 1824 2860 1832
rect 2842 1813 2846 1824
rect 2805 1801 2814 1813
rect 2725 1787 2734 1799
rect 2725 1771 2731 1787
rect 2703 1764 2717 1771
rect 2713 1744 2717 1764
rect 2723 1764 2731 1771
rect 2723 1744 2727 1764
rect 2785 1724 2789 1801
rect 2805 1724 2809 1801
rect 2842 1756 2846 1801
rect 2864 1779 2868 1836
rect 2886 1833 2890 1876
rect 2886 1821 2893 1833
rect 2866 1767 2875 1779
rect 2842 1749 2855 1756
rect 2851 1744 2855 1749
rect 2871 1744 2875 1767
rect 2891 1744 2895 1821
rect 2951 1793 2955 1876
rect 3113 1873 3117 1896
rect 3109 1866 3117 1873
rect 3109 1837 3113 1866
rect 3121 1856 3125 1896
rect 3141 1844 3145 1876
rect 3149 1872 3153 1876
rect 3149 1870 3185 1872
rect 3149 1868 3173 1870
rect 3037 1813 3041 1836
rect 3026 1801 3041 1813
rect 3045 1813 3049 1836
rect 3091 1824 3095 1836
rect 3109 1831 3117 1837
rect 3045 1801 3054 1813
rect 3091 1812 3093 1824
rect 2946 1781 2955 1793
rect 2951 1724 2955 1781
rect 3025 1724 3029 1801
rect 3045 1724 3049 1801
rect 3091 1744 3095 1812
rect 3113 1785 3117 1831
rect 3113 1724 3117 1773
rect 3141 1749 3147 1844
rect 3123 1745 3147 1749
rect 3123 1724 3127 1745
rect 3143 1740 3161 1741
rect 3143 1736 3173 1740
rect 3143 1724 3147 1736
rect 3181 1732 3185 1858
rect 3195 1850 3199 1876
rect 3215 1870 3219 1876
rect 3151 1728 3185 1732
rect 3151 1724 3155 1728
rect 3197 1724 3201 1838
rect 3213 1748 3217 1858
rect 3227 1836 3231 1876
rect 3222 1824 3225 1836
rect 3222 1760 3226 1824
rect 3247 1817 3251 1876
rect 3242 1809 3251 1817
rect 3242 1780 3246 1809
rect 3261 1794 3265 1876
rect 3281 1793 3285 1836
rect 3336 1832 3340 1836
rect 3322 1824 3340 1832
rect 3322 1813 3326 1824
rect 3222 1756 3255 1760
rect 3221 1736 3223 1748
rect 3219 1724 3223 1736
rect 3229 1736 3231 1748
rect 3229 1724 3233 1736
rect 3251 1724 3255 1756
rect 3261 1724 3265 1782
rect 3281 1744 3285 1781
rect 3322 1756 3326 1801
rect 3344 1779 3348 1836
rect 3366 1833 3370 1876
rect 3366 1821 3373 1833
rect 3346 1767 3355 1779
rect 3322 1749 3335 1756
rect 3331 1744 3335 1749
rect 3351 1744 3355 1767
rect 3371 1744 3375 1821
rect 3431 1799 3435 1876
rect 3426 1787 3435 1799
rect 3429 1771 3435 1787
rect 3451 1799 3455 1876
rect 3533 1873 3537 1896
rect 3529 1866 3537 1873
rect 3529 1837 3533 1866
rect 3541 1856 3545 1896
rect 3561 1844 3565 1876
rect 3569 1872 3573 1876
rect 3569 1870 3605 1872
rect 3569 1868 3593 1870
rect 3511 1824 3515 1836
rect 3529 1831 3537 1837
rect 3511 1812 3513 1824
rect 3451 1787 3454 1799
rect 3451 1771 3457 1787
rect 3429 1764 3437 1771
rect 3433 1744 3437 1764
rect 3443 1764 3457 1771
rect 3443 1744 3447 1764
rect 3511 1744 3515 1812
rect 3533 1785 3537 1831
rect 3533 1724 3537 1773
rect 3561 1749 3567 1844
rect 3543 1745 3567 1749
rect 3543 1724 3547 1745
rect 3563 1740 3581 1741
rect 3563 1736 3593 1740
rect 3563 1724 3567 1736
rect 3601 1732 3605 1858
rect 3615 1850 3619 1876
rect 3635 1870 3639 1876
rect 3571 1728 3605 1732
rect 3571 1724 3575 1728
rect 3617 1724 3621 1838
rect 3633 1748 3637 1858
rect 3647 1836 3651 1876
rect 3642 1824 3645 1836
rect 3642 1760 3646 1824
rect 3667 1817 3671 1876
rect 3662 1809 3671 1817
rect 3662 1780 3666 1809
rect 3681 1794 3685 1876
rect 3701 1793 3705 1836
rect 3751 1813 3755 1876
rect 3773 1830 3777 1836
rect 3775 1818 3777 1830
rect 3746 1801 3755 1813
rect 3642 1756 3675 1760
rect 3641 1736 3643 1748
rect 3639 1724 3643 1736
rect 3649 1736 3651 1748
rect 3649 1724 3653 1736
rect 3671 1724 3675 1756
rect 3681 1724 3685 1782
rect 3701 1744 3705 1781
rect 3751 1724 3755 1801
rect 3845 1799 3849 1876
rect 3846 1787 3849 1799
rect 3843 1771 3849 1787
rect 3865 1799 3869 1876
rect 3930 1833 3934 1876
rect 3927 1821 3934 1833
rect 3865 1787 3874 1799
rect 3865 1771 3871 1787
rect 3843 1764 3857 1771
rect 3775 1750 3777 1762
rect 3773 1744 3777 1750
rect 3853 1744 3857 1764
rect 3863 1764 3871 1771
rect 3863 1744 3867 1764
rect 3925 1744 3929 1821
rect 3952 1779 3956 1836
rect 3960 1832 3964 1836
rect 4030 1833 4034 1876
rect 3960 1824 3978 1832
rect 3974 1813 3978 1824
rect 4027 1821 4034 1833
rect 3945 1767 3954 1779
rect 3945 1744 3949 1767
rect 3974 1756 3978 1801
rect 3965 1749 3978 1756
rect 3965 1744 3969 1749
rect 4025 1744 4029 1821
rect 4052 1779 4056 1836
rect 4060 1832 4064 1836
rect 4111 1832 4115 1836
rect 4060 1824 4078 1832
rect 4074 1813 4078 1824
rect 4102 1827 4115 1832
rect 4045 1767 4054 1779
rect 4045 1744 4049 1767
rect 4074 1756 4078 1801
rect 4102 1793 4106 1827
rect 4121 1813 4125 1836
rect 4141 1831 4145 1836
rect 4065 1749 4078 1756
rect 4065 1744 4069 1749
rect 4102 1736 4106 1781
rect 4121 1737 4125 1801
rect 4225 1793 4229 1876
rect 4473 1873 4477 1896
rect 4469 1866 4477 1873
rect 4469 1837 4473 1866
rect 4481 1856 4485 1896
rect 4501 1844 4505 1876
rect 4509 1872 4513 1876
rect 4509 1870 4545 1872
rect 4509 1868 4533 1870
rect 4271 1822 4275 1836
rect 4291 1822 4295 1836
rect 4259 1816 4275 1822
rect 4280 1816 4295 1822
rect 4225 1781 4234 1793
rect 4145 1752 4155 1764
rect 4151 1744 4155 1752
rect 4102 1731 4115 1736
rect 4121 1731 4135 1737
rect 4111 1724 4115 1731
rect 4131 1724 4135 1731
rect 4225 1724 4229 1781
rect 4259 1779 4266 1816
rect 4280 1793 4286 1816
rect 4259 1754 4266 1767
rect 4259 1748 4278 1754
rect 4274 1744 4278 1748
rect 4282 1744 4286 1781
rect 4311 1779 4315 1836
rect 4397 1813 4401 1836
rect 4386 1801 4401 1813
rect 4405 1813 4409 1836
rect 4451 1824 4455 1836
rect 4469 1831 4477 1837
rect 4405 1801 4414 1813
rect 4451 1812 4453 1824
rect 4306 1767 4315 1779
rect 4304 1724 4308 1767
rect 4385 1724 4389 1801
rect 4405 1724 4409 1801
rect 4451 1744 4455 1812
rect 4473 1785 4477 1831
rect 4473 1724 4477 1773
rect 4501 1749 4507 1844
rect 4483 1745 4507 1749
rect 4483 1724 4487 1745
rect 4503 1740 4521 1741
rect 4503 1736 4533 1740
rect 4503 1724 4507 1736
rect 4541 1732 4545 1858
rect 4555 1850 4559 1876
rect 4575 1870 4579 1876
rect 4511 1728 4545 1732
rect 4511 1724 4515 1728
rect 4557 1724 4561 1838
rect 4573 1748 4577 1858
rect 4587 1836 4591 1876
rect 4582 1824 4585 1836
rect 4582 1760 4586 1824
rect 4607 1817 4611 1876
rect 4602 1809 4611 1817
rect 4602 1780 4606 1809
rect 4621 1794 4625 1876
rect 4641 1793 4645 1836
rect 4705 1799 4709 1876
rect 4582 1756 4615 1760
rect 4581 1736 4583 1748
rect 4579 1724 4583 1736
rect 4589 1736 4591 1748
rect 4589 1724 4593 1736
rect 4611 1724 4615 1756
rect 4621 1724 4625 1782
rect 4706 1787 4709 1799
rect 4641 1744 4645 1781
rect 4703 1771 4709 1787
rect 4725 1799 4729 1876
rect 4725 1787 4734 1799
rect 4725 1771 4731 1787
rect 4703 1764 4717 1771
rect 4713 1744 4717 1764
rect 4723 1764 4731 1771
rect 4723 1744 4727 1764
rect 66 1700 70 1704
rect 74 1700 78 1704
rect 94 1700 98 1704
rect 102 1700 106 1704
rect 151 1700 155 1704
rect 171 1700 175 1704
rect 191 1700 195 1704
rect 253 1700 257 1704
rect 263 1700 267 1704
rect 368 1700 372 1704
rect 376 1700 380 1704
rect 384 1700 388 1704
rect 434 1700 438 1704
rect 442 1700 446 1704
rect 462 1700 466 1704
rect 470 1700 474 1704
rect 551 1700 555 1704
rect 561 1700 565 1704
rect 581 1700 585 1704
rect 665 1700 669 1704
rect 711 1700 715 1704
rect 733 1700 737 1704
rect 805 1700 809 1704
rect 825 1700 829 1704
rect 845 1700 849 1704
rect 891 1700 895 1704
rect 911 1700 915 1704
rect 931 1700 935 1704
rect 992 1700 996 1704
rect 1000 1700 1004 1704
rect 1008 1700 1012 1704
rect 1091 1700 1095 1704
rect 1152 1700 1156 1704
rect 1160 1700 1164 1704
rect 1168 1700 1172 1704
rect 1252 1700 1256 1704
rect 1260 1700 1264 1704
rect 1268 1700 1272 1704
rect 1365 1700 1369 1704
rect 1446 1700 1450 1704
rect 1454 1700 1458 1704
rect 1474 1700 1478 1704
rect 1482 1700 1486 1704
rect 1532 1700 1536 1704
rect 1540 1700 1544 1704
rect 1548 1700 1552 1704
rect 1631 1700 1635 1704
rect 1705 1700 1709 1704
rect 1788 1700 1792 1704
rect 1796 1700 1800 1704
rect 1804 1700 1808 1704
rect 1851 1700 1855 1704
rect 1861 1700 1865 1704
rect 1881 1700 1885 1704
rect 1955 1700 1959 1704
rect 1975 1700 1979 1704
rect 1985 1700 1989 1704
rect 2007 1700 2011 1704
rect 2017 1700 2021 1704
rect 2039 1700 2043 1704
rect 2085 1700 2089 1704
rect 2093 1700 2097 1704
rect 2113 1700 2117 1704
rect 2123 1700 2127 1704
rect 2145 1700 2149 1704
rect 2205 1700 2209 1704
rect 2225 1700 2229 1704
rect 2271 1700 2275 1704
rect 2331 1700 2335 1704
rect 2351 1700 2355 1704
rect 2371 1700 2375 1704
rect 2431 1700 2435 1704
rect 2451 1700 2455 1704
rect 2511 1700 2515 1704
rect 2531 1700 2535 1704
rect 2591 1700 2595 1704
rect 2611 1700 2615 1704
rect 2631 1700 2635 1704
rect 2713 1700 2717 1704
rect 2723 1700 2727 1704
rect 2785 1700 2789 1704
rect 2805 1700 2809 1704
rect 2851 1700 2855 1704
rect 2871 1700 2875 1704
rect 2891 1700 2895 1704
rect 2951 1700 2955 1704
rect 3025 1700 3029 1704
rect 3045 1700 3049 1704
rect 3091 1700 3095 1704
rect 3113 1700 3117 1704
rect 3123 1700 3127 1704
rect 3143 1700 3147 1704
rect 3151 1700 3155 1704
rect 3197 1700 3201 1704
rect 3219 1700 3223 1704
rect 3229 1700 3233 1704
rect 3251 1700 3255 1704
rect 3261 1700 3265 1704
rect 3281 1700 3285 1704
rect 3331 1700 3335 1704
rect 3351 1700 3355 1704
rect 3371 1700 3375 1704
rect 3433 1700 3437 1704
rect 3443 1700 3447 1704
rect 3511 1700 3515 1704
rect 3533 1700 3537 1704
rect 3543 1700 3547 1704
rect 3563 1700 3567 1704
rect 3571 1700 3575 1704
rect 3617 1700 3621 1704
rect 3639 1700 3643 1704
rect 3649 1700 3653 1704
rect 3671 1700 3675 1704
rect 3681 1700 3685 1704
rect 3701 1700 3705 1704
rect 3751 1700 3755 1704
rect 3773 1700 3777 1704
rect 3853 1700 3857 1704
rect 3863 1700 3867 1704
rect 3925 1700 3929 1704
rect 3945 1700 3949 1704
rect 3965 1700 3969 1704
rect 4025 1700 4029 1704
rect 4045 1700 4049 1704
rect 4065 1700 4069 1704
rect 4111 1700 4115 1704
rect 4131 1700 4135 1704
rect 4151 1700 4155 1704
rect 4225 1700 4229 1704
rect 4274 1700 4278 1704
rect 4282 1700 4286 1704
rect 4304 1700 4308 1704
rect 4385 1700 4389 1704
rect 4405 1700 4409 1704
rect 4451 1700 4455 1704
rect 4473 1700 4477 1704
rect 4483 1700 4487 1704
rect 4503 1700 4507 1704
rect 4511 1700 4515 1704
rect 4557 1700 4561 1704
rect 4579 1700 4583 1704
rect 4589 1700 4593 1704
rect 4611 1700 4615 1704
rect 4621 1700 4625 1704
rect 4641 1700 4645 1704
rect 4713 1700 4717 1704
rect 4723 1700 4727 1704
rect 45 1676 49 1680
rect 112 1676 116 1680
rect 134 1676 138 1680
rect 142 1676 146 1680
rect 192 1676 196 1680
rect 200 1676 204 1680
rect 208 1676 212 1680
rect 293 1676 297 1680
rect 303 1676 307 1680
rect 385 1676 389 1680
rect 405 1676 409 1680
rect 425 1676 429 1680
rect 483 1676 487 1680
rect 505 1676 509 1680
rect 565 1676 569 1680
rect 612 1676 616 1680
rect 620 1676 624 1680
rect 628 1676 632 1680
rect 714 1676 718 1680
rect 722 1676 726 1680
rect 744 1676 748 1680
rect 812 1676 816 1680
rect 820 1676 824 1680
rect 828 1676 832 1680
rect 914 1676 918 1680
rect 922 1676 926 1680
rect 944 1676 948 1680
rect 1012 1676 1016 1680
rect 1020 1676 1024 1680
rect 1028 1676 1032 1680
rect 1125 1676 1129 1680
rect 1145 1676 1149 1680
rect 1165 1676 1169 1680
rect 1212 1676 1216 1680
rect 1220 1676 1224 1680
rect 1228 1676 1232 1680
rect 1314 1676 1318 1680
rect 1322 1676 1326 1680
rect 1344 1676 1348 1680
rect 1425 1676 1429 1680
rect 1472 1676 1476 1680
rect 1480 1676 1484 1680
rect 1488 1676 1492 1680
rect 1574 1676 1578 1680
rect 1582 1676 1586 1680
rect 1604 1676 1608 1680
rect 1672 1676 1676 1680
rect 1680 1676 1684 1680
rect 1688 1676 1692 1680
rect 1771 1676 1775 1680
rect 1791 1676 1795 1680
rect 1811 1676 1815 1680
rect 1892 1676 1896 1680
rect 1914 1676 1918 1680
rect 1922 1676 1926 1680
rect 1971 1676 1975 1680
rect 2032 1676 2036 1680
rect 2040 1676 2044 1680
rect 2048 1676 2052 1680
rect 2145 1676 2149 1680
rect 2165 1676 2169 1680
rect 2185 1676 2189 1680
rect 2231 1676 2235 1680
rect 2291 1676 2295 1680
rect 2313 1676 2317 1680
rect 2323 1676 2327 1680
rect 2343 1676 2347 1680
rect 2351 1676 2355 1680
rect 2397 1676 2401 1680
rect 2419 1676 2423 1680
rect 2429 1676 2433 1680
rect 2451 1676 2455 1680
rect 2461 1676 2465 1680
rect 2481 1676 2485 1680
rect 2545 1676 2549 1680
rect 2565 1676 2569 1680
rect 2585 1676 2589 1680
rect 2655 1676 2659 1680
rect 2675 1676 2679 1680
rect 2685 1676 2689 1680
rect 2731 1676 2735 1680
rect 2751 1676 2755 1680
rect 2814 1676 2818 1680
rect 2822 1676 2826 1680
rect 2844 1676 2848 1680
rect 2925 1676 2929 1680
rect 2945 1676 2949 1680
rect 3005 1676 3009 1680
rect 3065 1676 3069 1680
rect 3111 1676 3115 1680
rect 3131 1676 3135 1680
rect 3151 1676 3155 1680
rect 3213 1676 3217 1680
rect 3223 1676 3227 1680
rect 3313 1676 3317 1680
rect 3323 1676 3327 1680
rect 3385 1676 3389 1680
rect 3405 1676 3409 1680
rect 3425 1676 3429 1680
rect 3475 1676 3479 1680
rect 3495 1676 3499 1680
rect 3505 1676 3509 1680
rect 3527 1676 3531 1680
rect 3537 1676 3541 1680
rect 3559 1676 3563 1680
rect 3605 1676 3609 1680
rect 3613 1676 3617 1680
rect 3633 1676 3637 1680
rect 3643 1676 3647 1680
rect 3665 1676 3669 1680
rect 3711 1676 3715 1680
rect 3785 1676 3789 1680
rect 3845 1676 3849 1680
rect 3865 1676 3869 1680
rect 3885 1676 3889 1680
rect 3931 1676 3935 1680
rect 3951 1676 3955 1680
rect 4011 1676 4015 1680
rect 4031 1676 4035 1680
rect 4091 1676 4095 1680
rect 4154 1676 4158 1680
rect 4162 1676 4166 1680
rect 4184 1676 4188 1680
rect 4251 1676 4255 1680
rect 4271 1676 4275 1680
rect 4334 1676 4338 1680
rect 4342 1676 4346 1680
rect 4364 1676 4368 1680
rect 4431 1676 4435 1680
rect 4491 1676 4495 1680
rect 4565 1676 4569 1680
rect 4611 1676 4615 1680
rect 4631 1676 4635 1680
rect 4651 1676 4655 1680
rect 4713 1676 4717 1680
rect 4723 1676 4727 1680
rect 45 1599 49 1656
rect 112 1613 116 1656
rect 105 1601 114 1613
rect 45 1587 54 1599
rect 45 1504 49 1587
rect 105 1544 109 1601
rect 134 1599 138 1636
rect 142 1632 146 1636
rect 142 1626 161 1632
rect 154 1613 161 1626
rect 293 1616 297 1636
rect 134 1564 140 1587
rect 154 1564 161 1601
rect 125 1558 140 1564
rect 145 1558 161 1564
rect 192 1559 196 1616
rect 125 1544 129 1558
rect 145 1544 149 1558
rect 186 1547 196 1559
rect 180 1516 186 1547
rect 200 1539 204 1616
rect 208 1559 212 1616
rect 289 1609 297 1616
rect 303 1616 307 1636
rect 303 1609 317 1616
rect 289 1593 295 1609
rect 286 1581 295 1593
rect 208 1547 215 1559
rect 227 1547 235 1559
rect 200 1520 206 1527
rect 200 1516 215 1520
rect 180 1512 195 1516
rect 191 1504 195 1512
rect 211 1504 215 1516
rect 231 1504 235 1547
rect 291 1504 295 1581
rect 311 1593 317 1609
rect 311 1581 314 1593
rect 311 1504 315 1581
rect 385 1559 389 1636
rect 405 1613 409 1636
rect 425 1631 429 1636
rect 425 1624 438 1631
rect 405 1601 414 1613
rect 387 1547 394 1559
rect 390 1504 394 1547
rect 412 1544 416 1601
rect 434 1579 438 1624
rect 483 1630 487 1636
rect 483 1618 485 1630
rect 505 1579 509 1656
rect 565 1599 569 1656
rect 714 1632 718 1636
rect 699 1626 718 1632
rect 565 1587 574 1599
rect 505 1567 514 1579
rect 434 1556 438 1567
rect 420 1548 438 1556
rect 483 1550 485 1562
rect 420 1544 424 1548
rect 483 1544 487 1550
rect 505 1504 509 1567
rect 565 1504 569 1587
rect 612 1559 616 1616
rect 606 1547 616 1559
rect 600 1516 606 1547
rect 620 1539 624 1616
rect 628 1559 632 1616
rect 699 1613 706 1626
rect 699 1564 706 1601
rect 722 1599 726 1636
rect 744 1613 748 1656
rect 914 1632 918 1636
rect 899 1626 918 1632
rect 746 1601 755 1613
rect 720 1564 726 1587
rect 628 1547 635 1559
rect 647 1547 655 1559
rect 699 1558 715 1564
rect 720 1558 735 1564
rect 620 1520 626 1527
rect 620 1516 635 1520
rect 600 1512 615 1516
rect 611 1504 615 1512
rect 631 1504 635 1516
rect 651 1504 655 1547
rect 711 1544 715 1558
rect 731 1544 735 1558
rect 751 1544 755 1601
rect 812 1559 816 1616
rect 806 1547 816 1559
rect 800 1516 806 1547
rect 820 1539 824 1616
rect 828 1559 832 1616
rect 899 1613 906 1626
rect 899 1564 906 1601
rect 922 1599 926 1636
rect 944 1613 948 1656
rect 946 1601 955 1613
rect 920 1564 926 1587
rect 828 1547 835 1559
rect 847 1547 855 1559
rect 899 1558 915 1564
rect 920 1558 935 1564
rect 820 1520 826 1527
rect 820 1516 835 1520
rect 800 1512 815 1516
rect 811 1504 815 1512
rect 831 1504 835 1516
rect 851 1504 855 1547
rect 911 1544 915 1558
rect 931 1544 935 1558
rect 951 1544 955 1601
rect 1012 1559 1016 1616
rect 1006 1547 1016 1559
rect 1000 1516 1006 1547
rect 1020 1539 1024 1616
rect 1028 1559 1032 1616
rect 1125 1559 1129 1636
rect 1145 1613 1149 1636
rect 1165 1631 1169 1636
rect 1165 1624 1178 1631
rect 1145 1601 1154 1613
rect 1028 1547 1035 1559
rect 1047 1547 1055 1559
rect 1127 1547 1134 1559
rect 1020 1520 1026 1527
rect 1020 1516 1035 1520
rect 1000 1512 1015 1516
rect 1011 1504 1015 1512
rect 1031 1504 1035 1516
rect 1051 1504 1055 1547
rect 1130 1504 1134 1547
rect 1152 1544 1156 1601
rect 1174 1579 1178 1624
rect 1314 1632 1318 1636
rect 1299 1626 1318 1632
rect 1174 1556 1178 1567
rect 1212 1559 1216 1616
rect 1160 1548 1178 1556
rect 1160 1544 1164 1548
rect 1206 1547 1216 1559
rect 1200 1516 1206 1547
rect 1220 1539 1224 1616
rect 1228 1559 1232 1616
rect 1299 1613 1306 1626
rect 1299 1564 1306 1601
rect 1322 1599 1326 1636
rect 1344 1613 1348 1656
rect 1346 1601 1355 1613
rect 1320 1564 1326 1587
rect 1228 1547 1235 1559
rect 1247 1547 1255 1559
rect 1299 1558 1315 1564
rect 1320 1558 1335 1564
rect 1220 1520 1226 1527
rect 1220 1516 1235 1520
rect 1200 1512 1215 1516
rect 1211 1504 1215 1512
rect 1231 1504 1235 1516
rect 1251 1504 1255 1547
rect 1311 1544 1315 1558
rect 1331 1544 1335 1558
rect 1351 1544 1355 1601
rect 1425 1599 1429 1656
rect 1574 1632 1578 1636
rect 1559 1626 1578 1632
rect 1425 1587 1434 1599
rect 1425 1504 1429 1587
rect 1472 1559 1476 1616
rect 1466 1547 1476 1559
rect 1460 1516 1466 1547
rect 1480 1539 1484 1616
rect 1488 1559 1492 1616
rect 1559 1613 1566 1626
rect 1559 1564 1566 1601
rect 1582 1599 1586 1636
rect 1604 1613 1608 1656
rect 1771 1631 1775 1636
rect 1762 1624 1775 1631
rect 1606 1601 1615 1613
rect 1580 1564 1586 1587
rect 1488 1547 1495 1559
rect 1507 1547 1515 1559
rect 1559 1558 1575 1564
rect 1580 1558 1595 1564
rect 1480 1520 1486 1527
rect 1480 1516 1495 1520
rect 1460 1512 1475 1516
rect 1471 1504 1475 1512
rect 1491 1504 1495 1516
rect 1511 1504 1515 1547
rect 1571 1544 1575 1558
rect 1591 1544 1595 1558
rect 1611 1544 1615 1601
rect 1672 1559 1676 1616
rect 1666 1547 1676 1559
rect 1660 1516 1666 1547
rect 1680 1539 1684 1616
rect 1688 1559 1692 1616
rect 1762 1579 1766 1624
rect 1791 1613 1795 1636
rect 1786 1601 1795 1613
rect 1688 1547 1695 1559
rect 1707 1547 1715 1559
rect 1762 1556 1766 1567
rect 1762 1548 1780 1556
rect 1680 1520 1686 1527
rect 1680 1516 1695 1520
rect 1660 1512 1675 1516
rect 1671 1504 1675 1512
rect 1691 1504 1695 1516
rect 1711 1504 1715 1547
rect 1776 1544 1780 1548
rect 1784 1544 1788 1601
rect 1811 1559 1815 1636
rect 1892 1613 1896 1656
rect 1885 1601 1894 1613
rect 1806 1547 1813 1559
rect 1806 1504 1810 1547
rect 1885 1544 1889 1601
rect 1914 1599 1918 1636
rect 1922 1632 1926 1636
rect 1922 1626 1941 1632
rect 1934 1613 1941 1626
rect 1914 1564 1920 1587
rect 1934 1564 1941 1601
rect 1971 1599 1975 1656
rect 1966 1587 1975 1599
rect 1905 1558 1920 1564
rect 1925 1558 1941 1564
rect 1905 1544 1909 1558
rect 1925 1544 1929 1558
rect 1971 1504 1975 1587
rect 2032 1559 2036 1616
rect 2026 1547 2036 1559
rect 2020 1516 2026 1547
rect 2040 1539 2044 1616
rect 2048 1559 2052 1616
rect 2145 1559 2149 1636
rect 2165 1613 2169 1636
rect 2185 1631 2189 1636
rect 2185 1624 2198 1631
rect 2165 1601 2174 1613
rect 2048 1547 2055 1559
rect 2067 1547 2075 1559
rect 2147 1547 2154 1559
rect 2040 1520 2046 1527
rect 2040 1516 2055 1520
rect 2020 1512 2035 1516
rect 2031 1504 2035 1512
rect 2051 1504 2055 1516
rect 2071 1504 2075 1547
rect 2150 1504 2154 1547
rect 2172 1544 2176 1601
rect 2194 1579 2198 1624
rect 2231 1599 2235 1656
rect 2226 1587 2235 1599
rect 2194 1556 2198 1567
rect 2180 1548 2198 1556
rect 2180 1544 2184 1548
rect 2231 1504 2235 1587
rect 2291 1568 2295 1636
rect 2313 1607 2317 1656
rect 2323 1635 2327 1656
rect 2343 1644 2347 1656
rect 2351 1652 2355 1656
rect 2351 1648 2385 1652
rect 2343 1640 2373 1644
rect 2343 1639 2361 1640
rect 2323 1631 2347 1635
rect 2291 1556 2293 1568
rect 2291 1544 2295 1556
rect 2313 1549 2317 1595
rect 2309 1543 2317 1549
rect 2309 1514 2313 1543
rect 2341 1536 2347 1631
rect 2309 1507 2317 1514
rect 2313 1484 2317 1507
rect 2321 1484 2325 1524
rect 2341 1504 2345 1536
rect 2381 1522 2385 1648
rect 2397 1542 2401 1656
rect 2419 1644 2423 1656
rect 2421 1632 2423 1644
rect 2429 1644 2433 1656
rect 2429 1632 2431 1644
rect 2349 1510 2373 1512
rect 2349 1508 2385 1510
rect 2349 1504 2353 1508
rect 2395 1504 2399 1530
rect 2413 1522 2417 1632
rect 2451 1624 2455 1656
rect 2422 1620 2455 1624
rect 2422 1556 2426 1620
rect 2442 1571 2446 1600
rect 2461 1598 2465 1656
rect 2481 1599 2485 1636
rect 2442 1563 2451 1571
rect 2422 1544 2425 1556
rect 2415 1504 2419 1510
rect 2427 1504 2431 1544
rect 2447 1504 2451 1563
rect 2461 1504 2465 1586
rect 2481 1544 2485 1587
rect 2545 1559 2549 1636
rect 2565 1613 2569 1636
rect 2585 1631 2589 1636
rect 2585 1624 2598 1631
rect 2655 1630 2659 1636
rect 2565 1601 2574 1613
rect 2547 1547 2554 1559
rect 2550 1504 2554 1547
rect 2572 1544 2576 1601
rect 2594 1579 2598 1624
rect 2641 1618 2653 1630
rect 2594 1556 2598 1567
rect 2580 1548 2598 1556
rect 2580 1544 2584 1548
rect 2641 1544 2645 1618
rect 2675 1593 2679 1636
rect 2666 1581 2679 1593
rect 2663 1504 2667 1581
rect 2685 1579 2689 1636
rect 2731 1579 2735 1656
rect 2751 1579 2755 1656
rect 2814 1632 2818 1636
rect 2799 1626 2818 1632
rect 2799 1613 2806 1626
rect 2685 1567 2694 1579
rect 2726 1567 2735 1579
rect 2685 1504 2689 1567
rect 2731 1544 2735 1567
rect 2739 1567 2754 1579
rect 2739 1544 2743 1567
rect 2799 1564 2806 1601
rect 2822 1599 2826 1636
rect 2844 1613 2848 1656
rect 2846 1601 2855 1613
rect 2820 1564 2826 1587
rect 2799 1558 2815 1564
rect 2820 1558 2835 1564
rect 2811 1544 2815 1558
rect 2831 1544 2835 1558
rect 2851 1544 2855 1601
rect 2925 1579 2929 1656
rect 2945 1579 2949 1656
rect 3005 1599 3009 1656
rect 3065 1599 3069 1656
rect 3111 1631 3115 1636
rect 3102 1624 3115 1631
rect 3005 1587 3014 1599
rect 3065 1587 3074 1599
rect 2926 1567 2941 1579
rect 2937 1544 2941 1567
rect 2945 1567 2954 1579
rect 2945 1544 2949 1567
rect 3005 1504 3009 1587
rect 3065 1504 3069 1587
rect 3102 1579 3106 1624
rect 3131 1613 3135 1636
rect 3126 1601 3135 1613
rect 3102 1556 3106 1567
rect 3102 1548 3120 1556
rect 3116 1544 3120 1548
rect 3124 1544 3128 1601
rect 3151 1559 3155 1636
rect 3213 1616 3217 1636
rect 3209 1609 3217 1616
rect 3223 1616 3227 1636
rect 3313 1616 3317 1636
rect 3223 1609 3237 1616
rect 3209 1593 3215 1609
rect 3206 1581 3215 1593
rect 3146 1547 3153 1559
rect 3146 1504 3150 1547
rect 3211 1504 3215 1581
rect 3231 1593 3237 1609
rect 3303 1609 3317 1616
rect 3323 1616 3327 1636
rect 3323 1609 3331 1616
rect 3303 1593 3309 1609
rect 3231 1581 3234 1593
rect 3306 1581 3309 1593
rect 3231 1504 3235 1581
rect 3305 1504 3309 1581
rect 3325 1593 3331 1609
rect 3325 1581 3334 1593
rect 3325 1504 3329 1581
rect 3385 1559 3389 1636
rect 3405 1613 3409 1636
rect 3425 1631 3429 1636
rect 3425 1624 3438 1631
rect 3405 1601 3414 1613
rect 3387 1547 3394 1559
rect 3390 1504 3394 1547
rect 3412 1544 3416 1601
rect 3434 1579 3438 1624
rect 3475 1599 3479 1636
rect 3495 1598 3499 1656
rect 3505 1624 3509 1656
rect 3527 1644 3531 1656
rect 3529 1632 3531 1644
rect 3537 1644 3541 1656
rect 3537 1632 3539 1644
rect 3505 1620 3538 1624
rect 3434 1556 3438 1567
rect 3420 1548 3438 1556
rect 3420 1544 3424 1548
rect 3475 1544 3479 1587
rect 3495 1504 3499 1586
rect 3514 1571 3518 1600
rect 3509 1563 3518 1571
rect 3509 1504 3513 1563
rect 3534 1556 3538 1620
rect 3535 1544 3538 1556
rect 3529 1504 3533 1544
rect 3543 1522 3547 1632
rect 3559 1542 3563 1656
rect 3605 1652 3609 1656
rect 3575 1648 3609 1652
rect 3541 1504 3545 1510
rect 3561 1504 3565 1530
rect 3575 1522 3579 1648
rect 3613 1644 3617 1656
rect 3587 1640 3617 1644
rect 3599 1639 3617 1640
rect 3633 1635 3637 1656
rect 3613 1631 3637 1635
rect 3613 1536 3619 1631
rect 3643 1607 3647 1656
rect 3643 1549 3647 1595
rect 3665 1568 3669 1636
rect 3711 1599 3715 1656
rect 3706 1587 3715 1599
rect 3667 1556 3669 1568
rect 3643 1543 3651 1549
rect 3665 1544 3669 1556
rect 3587 1510 3611 1512
rect 3575 1508 3611 1510
rect 3607 1504 3611 1508
rect 3615 1504 3619 1536
rect 3635 1484 3639 1524
rect 3647 1514 3651 1543
rect 3643 1507 3651 1514
rect 3643 1484 3647 1507
rect 3711 1504 3715 1587
rect 3785 1599 3789 1656
rect 3785 1587 3794 1599
rect 3785 1504 3789 1587
rect 3845 1559 3849 1636
rect 3865 1613 3869 1636
rect 3885 1631 3889 1636
rect 3885 1624 3898 1631
rect 3865 1601 3874 1613
rect 3847 1547 3854 1559
rect 3850 1504 3854 1547
rect 3872 1544 3876 1601
rect 3894 1579 3898 1624
rect 3931 1579 3935 1656
rect 3951 1579 3955 1656
rect 4011 1579 4015 1656
rect 4031 1579 4035 1656
rect 4091 1599 4095 1656
rect 4154 1632 4158 1636
rect 4139 1626 4158 1632
rect 4139 1613 4146 1626
rect 4086 1587 4095 1599
rect 3926 1567 3935 1579
rect 3894 1556 3898 1567
rect 3880 1548 3898 1556
rect 3880 1544 3884 1548
rect 3931 1544 3935 1567
rect 3939 1567 3954 1579
rect 4006 1567 4015 1579
rect 3939 1544 3943 1567
rect 4011 1544 4015 1567
rect 4019 1567 4034 1579
rect 4019 1544 4023 1567
rect 4091 1504 4095 1587
rect 4139 1564 4146 1601
rect 4162 1599 4166 1636
rect 4184 1613 4188 1656
rect 4186 1601 4195 1613
rect 4160 1564 4166 1587
rect 4139 1558 4155 1564
rect 4160 1558 4175 1564
rect 4151 1544 4155 1558
rect 4171 1544 4175 1558
rect 4191 1544 4195 1601
rect 4251 1579 4255 1656
rect 4271 1579 4275 1656
rect 4334 1632 4338 1636
rect 4319 1626 4338 1632
rect 4319 1613 4326 1626
rect 4246 1567 4255 1579
rect 4251 1544 4255 1567
rect 4259 1567 4274 1579
rect 4259 1544 4263 1567
rect 4319 1564 4326 1601
rect 4342 1599 4346 1636
rect 4364 1613 4368 1656
rect 4366 1601 4375 1613
rect 4340 1564 4346 1587
rect 4319 1558 4335 1564
rect 4340 1558 4355 1564
rect 4331 1544 4335 1558
rect 4351 1544 4355 1558
rect 4371 1544 4375 1601
rect 4431 1599 4435 1656
rect 4491 1599 4495 1656
rect 4426 1587 4435 1599
rect 4486 1587 4495 1599
rect 4431 1504 4435 1587
rect 4491 1504 4495 1587
rect 4565 1599 4569 1656
rect 4611 1631 4615 1636
rect 4602 1624 4615 1631
rect 4565 1587 4574 1599
rect 4565 1504 4569 1587
rect 4602 1579 4606 1624
rect 4631 1613 4635 1636
rect 4626 1601 4635 1613
rect 4602 1556 4606 1567
rect 4602 1548 4620 1556
rect 4616 1544 4620 1548
rect 4624 1544 4628 1601
rect 4651 1559 4655 1636
rect 4713 1616 4717 1636
rect 4709 1609 4717 1616
rect 4723 1616 4727 1636
rect 4723 1609 4737 1616
rect 4709 1593 4715 1609
rect 4706 1581 4715 1593
rect 4646 1547 4653 1559
rect 4646 1504 4650 1547
rect 4711 1504 4715 1581
rect 4731 1593 4737 1609
rect 4731 1581 4734 1593
rect 4731 1504 4735 1581
rect 45 1460 49 1464
rect 105 1460 109 1464
rect 125 1460 129 1464
rect 145 1460 149 1464
rect 191 1460 195 1464
rect 211 1460 215 1464
rect 231 1460 235 1464
rect 291 1460 295 1464
rect 311 1460 315 1464
rect 390 1460 394 1464
rect 412 1460 416 1464
rect 420 1460 424 1464
rect 483 1460 487 1464
rect 505 1460 509 1464
rect 565 1460 569 1464
rect 611 1460 615 1464
rect 631 1460 635 1464
rect 651 1460 655 1464
rect 711 1460 715 1464
rect 731 1460 735 1464
rect 751 1460 755 1464
rect 811 1460 815 1464
rect 831 1460 835 1464
rect 851 1460 855 1464
rect 911 1460 915 1464
rect 931 1460 935 1464
rect 951 1460 955 1464
rect 1011 1460 1015 1464
rect 1031 1460 1035 1464
rect 1051 1460 1055 1464
rect 1130 1460 1134 1464
rect 1152 1460 1156 1464
rect 1160 1460 1164 1464
rect 1211 1460 1215 1464
rect 1231 1460 1235 1464
rect 1251 1460 1255 1464
rect 1311 1460 1315 1464
rect 1331 1460 1335 1464
rect 1351 1460 1355 1464
rect 1425 1460 1429 1464
rect 1471 1460 1475 1464
rect 1491 1460 1495 1464
rect 1511 1460 1515 1464
rect 1571 1460 1575 1464
rect 1591 1460 1595 1464
rect 1611 1460 1615 1464
rect 1671 1460 1675 1464
rect 1691 1460 1695 1464
rect 1711 1460 1715 1464
rect 1776 1460 1780 1464
rect 1784 1460 1788 1464
rect 1806 1460 1810 1464
rect 1885 1460 1889 1464
rect 1905 1460 1909 1464
rect 1925 1460 1929 1464
rect 1971 1460 1975 1464
rect 2031 1460 2035 1464
rect 2051 1460 2055 1464
rect 2071 1460 2075 1464
rect 2150 1460 2154 1464
rect 2172 1460 2176 1464
rect 2180 1460 2184 1464
rect 2231 1460 2235 1464
rect 2291 1460 2295 1464
rect 2313 1460 2317 1464
rect 2321 1460 2325 1464
rect 2341 1460 2345 1464
rect 2349 1460 2353 1464
rect 2395 1460 2399 1464
rect 2415 1460 2419 1464
rect 2427 1460 2431 1464
rect 2447 1460 2451 1464
rect 2461 1460 2465 1464
rect 2481 1460 2485 1464
rect 2550 1460 2554 1464
rect 2572 1460 2576 1464
rect 2580 1460 2584 1464
rect 2641 1460 2645 1464
rect 2663 1460 2667 1464
rect 2685 1460 2689 1464
rect 2731 1460 2735 1464
rect 2739 1460 2743 1464
rect 2811 1460 2815 1464
rect 2831 1460 2835 1464
rect 2851 1460 2855 1464
rect 2937 1460 2941 1464
rect 2945 1460 2949 1464
rect 3005 1460 3009 1464
rect 3065 1460 3069 1464
rect 3116 1460 3120 1464
rect 3124 1460 3128 1464
rect 3146 1460 3150 1464
rect 3211 1460 3215 1464
rect 3231 1460 3235 1464
rect 3305 1460 3309 1464
rect 3325 1460 3329 1464
rect 3390 1460 3394 1464
rect 3412 1460 3416 1464
rect 3420 1460 3424 1464
rect 3475 1460 3479 1464
rect 3495 1460 3499 1464
rect 3509 1460 3513 1464
rect 3529 1460 3533 1464
rect 3541 1460 3545 1464
rect 3561 1460 3565 1464
rect 3607 1460 3611 1464
rect 3615 1460 3619 1464
rect 3635 1460 3639 1464
rect 3643 1460 3647 1464
rect 3665 1460 3669 1464
rect 3711 1460 3715 1464
rect 3785 1460 3789 1464
rect 3850 1460 3854 1464
rect 3872 1460 3876 1464
rect 3880 1460 3884 1464
rect 3931 1460 3935 1464
rect 3939 1460 3943 1464
rect 4011 1460 4015 1464
rect 4019 1460 4023 1464
rect 4091 1460 4095 1464
rect 4151 1460 4155 1464
rect 4171 1460 4175 1464
rect 4191 1460 4195 1464
rect 4251 1460 4255 1464
rect 4259 1460 4263 1464
rect 4331 1460 4335 1464
rect 4351 1460 4355 1464
rect 4371 1460 4375 1464
rect 4431 1460 4435 1464
rect 4491 1460 4495 1464
rect 4565 1460 4569 1464
rect 4616 1460 4620 1464
rect 4624 1460 4628 1464
rect 4646 1460 4650 1464
rect 4711 1460 4715 1464
rect 4731 1460 4735 1464
rect 45 1436 49 1440
rect 65 1436 69 1440
rect 85 1436 89 1440
rect 131 1436 135 1440
rect 151 1436 155 1440
rect 171 1436 175 1440
rect 231 1436 235 1440
rect 251 1436 255 1440
rect 271 1436 275 1440
rect 345 1436 349 1440
rect 365 1436 369 1440
rect 416 1436 420 1440
rect 424 1436 428 1440
rect 446 1436 450 1440
rect 511 1436 515 1440
rect 531 1436 535 1440
rect 551 1436 555 1440
rect 616 1436 620 1440
rect 624 1436 628 1440
rect 646 1436 650 1440
rect 716 1436 720 1440
rect 724 1436 728 1440
rect 746 1436 750 1440
rect 811 1436 815 1440
rect 833 1436 837 1440
rect 855 1436 859 1440
rect 925 1436 929 1440
rect 945 1436 949 1440
rect 991 1436 995 1440
rect 1011 1436 1015 1440
rect 1085 1436 1089 1440
rect 1105 1436 1109 1440
rect 1125 1436 1129 1440
rect 1185 1436 1189 1440
rect 1241 1436 1245 1440
rect 1263 1436 1267 1440
rect 1285 1436 1289 1440
rect 1336 1436 1340 1440
rect 1344 1436 1348 1440
rect 1366 1436 1370 1440
rect 1450 1436 1454 1440
rect 1472 1436 1476 1440
rect 1480 1436 1484 1440
rect 1531 1436 1535 1440
rect 1551 1436 1555 1440
rect 1616 1436 1620 1440
rect 1624 1436 1628 1440
rect 1646 1436 1650 1440
rect 1711 1436 1715 1440
rect 1731 1436 1735 1440
rect 1791 1436 1795 1440
rect 1811 1436 1815 1440
rect 1831 1436 1835 1440
rect 1891 1436 1895 1440
rect 1911 1436 1915 1440
rect 1931 1436 1935 1440
rect 1996 1436 2000 1440
rect 2004 1436 2008 1440
rect 2026 1436 2030 1440
rect 2091 1436 2095 1440
rect 2151 1436 2155 1440
rect 2171 1436 2175 1440
rect 2191 1436 2195 1440
rect 2251 1436 2255 1440
rect 2271 1436 2275 1440
rect 2331 1436 2335 1440
rect 2341 1436 2345 1440
rect 2361 1436 2365 1440
rect 2445 1436 2449 1440
rect 2465 1436 2469 1440
rect 2511 1436 2515 1440
rect 2583 1436 2587 1440
rect 2605 1436 2609 1440
rect 2656 1436 2660 1440
rect 2664 1436 2668 1440
rect 2686 1436 2690 1440
rect 2775 1436 2779 1440
rect 2785 1436 2789 1440
rect 2815 1436 2819 1440
rect 2825 1436 2829 1440
rect 2875 1436 2879 1440
rect 2895 1436 2899 1440
rect 2909 1436 2913 1440
rect 2929 1436 2933 1440
rect 2941 1436 2945 1440
rect 2961 1436 2965 1440
rect 3007 1436 3011 1440
rect 3015 1436 3019 1440
rect 3035 1436 3039 1440
rect 3043 1436 3047 1440
rect 3065 1436 3069 1440
rect 3137 1436 3141 1440
rect 3145 1436 3149 1440
rect 3205 1436 3209 1440
rect 3225 1436 3229 1440
rect 3245 1436 3249 1440
rect 3295 1436 3299 1440
rect 3315 1436 3319 1440
rect 3329 1436 3333 1440
rect 3349 1436 3353 1440
rect 3361 1436 3365 1440
rect 3381 1436 3385 1440
rect 3427 1436 3431 1440
rect 3435 1436 3439 1440
rect 3455 1436 3459 1440
rect 3463 1436 3467 1440
rect 3485 1436 3489 1440
rect 3545 1436 3549 1440
rect 3617 1436 3621 1440
rect 3625 1436 3629 1440
rect 3697 1436 3701 1440
rect 3705 1436 3709 1440
rect 3751 1436 3755 1440
rect 3811 1436 3815 1440
rect 3833 1436 3837 1440
rect 3841 1436 3845 1440
rect 3861 1436 3865 1440
rect 3869 1436 3873 1440
rect 3915 1436 3919 1440
rect 3935 1436 3939 1440
rect 3947 1436 3951 1440
rect 3967 1436 3971 1440
rect 3981 1436 3985 1440
rect 4001 1436 4005 1440
rect 4056 1436 4060 1440
rect 4064 1436 4068 1440
rect 4086 1436 4090 1440
rect 4151 1436 4155 1440
rect 4171 1436 4175 1440
rect 4243 1436 4247 1440
rect 4265 1436 4269 1440
rect 4325 1436 4329 1440
rect 4345 1436 4349 1440
rect 4410 1436 4414 1440
rect 4432 1436 4436 1440
rect 4440 1436 4444 1440
rect 4510 1436 4514 1440
rect 4532 1436 4536 1440
rect 4540 1436 4544 1440
rect 4591 1436 4595 1440
rect 4599 1436 4603 1440
rect 4671 1436 4675 1440
rect 4745 1436 4749 1440
rect 131 1388 135 1396
rect 120 1384 135 1388
rect 151 1384 155 1396
rect 45 1299 49 1356
rect 65 1342 69 1356
rect 85 1342 89 1356
rect 120 1353 126 1384
rect 140 1380 155 1384
rect 140 1373 146 1380
rect 65 1336 80 1342
rect 85 1336 101 1342
rect 126 1341 136 1353
rect 74 1313 80 1336
rect 45 1287 54 1299
rect 52 1244 56 1287
rect 74 1264 78 1301
rect 94 1299 101 1336
rect 94 1274 101 1287
rect 132 1284 136 1341
rect 140 1284 144 1361
rect 171 1353 175 1396
rect 231 1388 235 1396
rect 220 1384 235 1388
rect 251 1384 255 1396
rect 220 1353 226 1384
rect 240 1380 255 1384
rect 240 1373 246 1380
rect 148 1341 155 1353
rect 167 1341 175 1353
rect 226 1341 236 1353
rect 148 1284 152 1341
rect 232 1284 236 1341
rect 240 1284 244 1361
rect 271 1353 275 1396
rect 248 1341 255 1353
rect 267 1341 275 1353
rect 248 1284 252 1341
rect 345 1319 349 1396
rect 346 1307 349 1319
rect 343 1291 349 1307
rect 365 1319 369 1396
rect 416 1352 420 1356
rect 402 1344 420 1352
rect 402 1333 406 1344
rect 365 1307 374 1319
rect 365 1291 371 1307
rect 343 1284 357 1291
rect 82 1268 101 1274
rect 82 1264 86 1268
rect 353 1264 357 1284
rect 363 1284 371 1291
rect 363 1264 367 1284
rect 402 1276 406 1321
rect 424 1299 428 1356
rect 446 1353 450 1396
rect 446 1341 453 1353
rect 511 1342 515 1356
rect 531 1342 535 1356
rect 426 1287 435 1299
rect 402 1269 415 1276
rect 411 1264 415 1269
rect 431 1264 435 1287
rect 451 1264 455 1341
rect 499 1336 515 1342
rect 520 1336 535 1342
rect 499 1299 506 1336
rect 520 1313 526 1336
rect 499 1274 506 1287
rect 499 1268 518 1274
rect 514 1264 518 1268
rect 522 1264 526 1301
rect 551 1299 555 1356
rect 616 1352 620 1356
rect 602 1344 620 1352
rect 602 1333 606 1344
rect 546 1287 555 1299
rect 544 1244 548 1287
rect 602 1276 606 1321
rect 624 1299 628 1356
rect 646 1353 650 1396
rect 646 1341 653 1353
rect 716 1352 720 1356
rect 702 1344 720 1352
rect 626 1287 635 1299
rect 602 1269 615 1276
rect 611 1264 615 1269
rect 631 1264 635 1287
rect 651 1264 655 1341
rect 702 1333 706 1344
rect 702 1276 706 1321
rect 724 1299 728 1356
rect 746 1353 750 1396
rect 746 1341 753 1353
rect 726 1287 735 1299
rect 702 1269 715 1276
rect 711 1264 715 1269
rect 731 1264 735 1287
rect 751 1264 755 1341
rect 811 1333 815 1396
rect 806 1321 815 1333
rect 811 1264 815 1321
rect 833 1319 837 1396
rect 821 1307 834 1319
rect 821 1264 825 1307
rect 855 1282 859 1356
rect 925 1319 929 1396
rect 926 1307 929 1319
rect 923 1291 929 1307
rect 945 1319 949 1396
rect 991 1319 995 1396
rect 945 1307 954 1319
rect 986 1307 995 1319
rect 945 1291 951 1307
rect 923 1284 937 1291
rect 847 1270 859 1282
rect 841 1264 845 1270
rect 933 1264 937 1284
rect 943 1284 951 1291
rect 989 1291 995 1307
rect 1011 1319 1015 1396
rect 1085 1353 1089 1396
rect 1105 1384 1109 1396
rect 1125 1388 1129 1396
rect 1125 1384 1140 1388
rect 1105 1380 1120 1384
rect 1114 1373 1120 1380
rect 1085 1341 1093 1353
rect 1105 1341 1112 1353
rect 1011 1307 1014 1319
rect 1011 1291 1017 1307
rect 989 1284 997 1291
rect 943 1264 947 1284
rect 993 1264 997 1284
rect 1003 1284 1017 1291
rect 1108 1284 1112 1341
rect 1116 1284 1120 1361
rect 1134 1353 1140 1384
rect 1124 1341 1134 1353
rect 1124 1284 1128 1341
rect 1185 1313 1189 1396
rect 1185 1301 1194 1313
rect 1003 1264 1007 1284
rect 1185 1244 1189 1301
rect 1241 1282 1245 1356
rect 1263 1319 1267 1396
rect 1285 1333 1289 1396
rect 1336 1352 1340 1356
rect 1322 1344 1340 1352
rect 1322 1333 1326 1344
rect 1285 1321 1294 1333
rect 1266 1307 1279 1319
rect 1241 1270 1253 1282
rect 1255 1264 1259 1270
rect 1275 1264 1279 1307
rect 1285 1264 1289 1321
rect 1322 1276 1326 1321
rect 1344 1299 1348 1356
rect 1366 1353 1370 1396
rect 1450 1353 1454 1396
rect 1366 1341 1373 1353
rect 1447 1341 1454 1353
rect 1346 1287 1355 1299
rect 1322 1269 1335 1276
rect 1331 1264 1335 1269
rect 1351 1264 1355 1287
rect 1371 1264 1375 1341
rect 1445 1264 1449 1341
rect 1472 1299 1476 1356
rect 1480 1352 1484 1356
rect 1480 1344 1498 1352
rect 1494 1333 1498 1344
rect 1465 1287 1474 1299
rect 1465 1264 1469 1287
rect 1494 1276 1498 1321
rect 1531 1319 1535 1396
rect 1526 1307 1535 1319
rect 1529 1291 1535 1307
rect 1551 1319 1555 1396
rect 1616 1352 1620 1356
rect 1602 1344 1620 1352
rect 1602 1333 1606 1344
rect 1551 1307 1554 1319
rect 1551 1291 1557 1307
rect 1529 1284 1537 1291
rect 1485 1269 1498 1276
rect 1485 1264 1489 1269
rect 1533 1264 1537 1284
rect 1543 1284 1557 1291
rect 1543 1264 1547 1284
rect 1602 1276 1606 1321
rect 1624 1299 1628 1356
rect 1646 1353 1650 1396
rect 1646 1341 1653 1353
rect 1626 1287 1635 1299
rect 1602 1269 1615 1276
rect 1611 1264 1615 1269
rect 1631 1264 1635 1287
rect 1651 1264 1655 1341
rect 1711 1319 1715 1396
rect 1706 1307 1715 1319
rect 1709 1291 1715 1307
rect 1731 1319 1735 1396
rect 1891 1388 1895 1396
rect 1880 1384 1895 1388
rect 1911 1384 1915 1396
rect 1791 1342 1795 1356
rect 1811 1342 1815 1356
rect 1779 1336 1795 1342
rect 1800 1336 1815 1342
rect 1731 1307 1734 1319
rect 1731 1291 1737 1307
rect 1779 1299 1786 1336
rect 1800 1313 1806 1336
rect 1709 1284 1717 1291
rect 1713 1264 1717 1284
rect 1723 1284 1737 1291
rect 1723 1264 1727 1284
rect 1779 1274 1786 1287
rect 1779 1268 1798 1274
rect 1794 1264 1798 1268
rect 1802 1264 1806 1301
rect 1831 1299 1835 1356
rect 1880 1353 1886 1384
rect 1900 1380 1915 1384
rect 1900 1373 1906 1380
rect 1886 1341 1896 1353
rect 1826 1287 1835 1299
rect 1824 1244 1828 1287
rect 1892 1284 1896 1341
rect 1900 1284 1904 1361
rect 1931 1353 1935 1396
rect 1908 1341 1915 1353
rect 1927 1341 1935 1353
rect 1996 1352 2000 1356
rect 1982 1344 2000 1352
rect 1908 1284 1912 1341
rect 1982 1333 1986 1344
rect 1982 1276 1986 1321
rect 2004 1299 2008 1356
rect 2026 1353 2030 1396
rect 2026 1341 2033 1353
rect 2006 1287 2015 1299
rect 1982 1269 1995 1276
rect 1991 1264 1995 1269
rect 2011 1264 2015 1287
rect 2031 1264 2035 1341
rect 2091 1313 2095 1396
rect 2151 1388 2155 1396
rect 2140 1384 2155 1388
rect 2171 1384 2175 1396
rect 2140 1353 2146 1384
rect 2160 1380 2175 1384
rect 2160 1373 2166 1380
rect 2146 1341 2156 1353
rect 2086 1301 2095 1313
rect 2091 1244 2095 1301
rect 2152 1284 2156 1341
rect 2160 1284 2164 1361
rect 2191 1353 2195 1396
rect 2168 1341 2175 1353
rect 2187 1341 2195 1353
rect 2168 1284 2172 1341
rect 2251 1319 2255 1396
rect 2246 1307 2255 1319
rect 2249 1291 2255 1307
rect 2271 1319 2275 1396
rect 2331 1352 2335 1356
rect 2322 1347 2335 1352
rect 2271 1307 2274 1319
rect 2322 1313 2326 1347
rect 2341 1333 2345 1356
rect 2361 1351 2365 1356
rect 2271 1291 2277 1307
rect 2249 1284 2257 1291
rect 2253 1264 2257 1284
rect 2263 1284 2277 1291
rect 2263 1264 2267 1284
rect 2322 1256 2326 1301
rect 2341 1257 2345 1321
rect 2445 1319 2449 1396
rect 2446 1307 2449 1319
rect 2443 1291 2449 1307
rect 2465 1319 2469 1396
rect 2465 1307 2474 1319
rect 2511 1313 2515 1396
rect 2583 1350 2587 1356
rect 2583 1338 2585 1350
rect 2465 1291 2471 1307
rect 2506 1301 2515 1313
rect 2443 1284 2457 1291
rect 2365 1272 2375 1284
rect 2371 1264 2375 1272
rect 2453 1264 2457 1284
rect 2463 1284 2471 1291
rect 2463 1264 2467 1284
rect 2322 1251 2335 1256
rect 2341 1251 2355 1257
rect 2331 1244 2335 1251
rect 2351 1244 2355 1251
rect 2511 1244 2515 1301
rect 2605 1333 2609 1396
rect 2656 1352 2660 1356
rect 2642 1344 2660 1352
rect 2642 1333 2646 1344
rect 2605 1321 2614 1333
rect 2583 1270 2585 1282
rect 2583 1264 2587 1270
rect 2605 1244 2609 1321
rect 2642 1276 2646 1321
rect 2664 1299 2668 1356
rect 2686 1353 2690 1396
rect 2686 1341 2693 1353
rect 2775 1352 2779 1356
rect 2765 1348 2779 1352
rect 2666 1287 2675 1299
rect 2642 1269 2655 1276
rect 2651 1264 2655 1269
rect 2671 1264 2675 1287
rect 2691 1264 2695 1341
rect 2765 1333 2769 1348
rect 2767 1321 2769 1333
rect 2765 1264 2769 1321
rect 2785 1299 2789 1356
rect 2815 1352 2819 1356
rect 2805 1348 2819 1352
rect 2825 1352 2829 1356
rect 2825 1348 2839 1352
rect 2805 1299 2811 1348
rect 2834 1333 2839 1348
rect 2805 1287 2814 1299
rect 2785 1264 2789 1287
rect 2805 1264 2809 1287
rect 2834 1275 2840 1321
rect 2875 1313 2879 1356
rect 2895 1314 2899 1396
rect 2909 1337 2913 1396
rect 2929 1356 2933 1396
rect 2941 1390 2945 1396
rect 2935 1344 2938 1356
rect 2909 1329 2918 1337
rect 2825 1271 2840 1275
rect 2825 1264 2829 1271
rect 2875 1264 2879 1301
rect 2895 1244 2899 1302
rect 2914 1300 2918 1329
rect 2934 1280 2938 1344
rect 2905 1276 2938 1280
rect 2905 1244 2909 1276
rect 2943 1268 2947 1378
rect 2961 1370 2965 1396
rect 3007 1392 3011 1396
rect 2975 1390 3011 1392
rect 2987 1388 3011 1390
rect 2929 1256 2931 1268
rect 2927 1244 2931 1256
rect 2937 1256 2939 1268
rect 2937 1244 2941 1256
rect 2959 1244 2963 1358
rect 2975 1252 2979 1378
rect 3015 1364 3019 1396
rect 3035 1376 3039 1416
rect 3043 1393 3047 1416
rect 3043 1386 3051 1393
rect 3013 1269 3019 1364
rect 3047 1357 3051 1386
rect 3043 1351 3051 1357
rect 3043 1305 3047 1351
rect 3065 1344 3069 1356
rect 3067 1332 3069 1344
rect 3137 1333 3141 1356
rect 3013 1265 3037 1269
rect 2999 1260 3017 1261
rect 2987 1256 3017 1260
rect 2975 1248 3009 1252
rect 3005 1244 3009 1248
rect 3013 1244 3017 1256
rect 3033 1244 3037 1265
rect 3043 1244 3047 1293
rect 3065 1264 3069 1332
rect 3126 1321 3141 1333
rect 3145 1333 3149 1356
rect 3145 1321 3154 1333
rect 3125 1244 3129 1321
rect 3145 1244 3149 1321
rect 3205 1299 3209 1356
rect 3225 1342 3229 1356
rect 3245 1342 3249 1356
rect 3225 1336 3240 1342
rect 3245 1336 3261 1342
rect 3234 1313 3240 1336
rect 3205 1287 3214 1299
rect 3212 1244 3216 1287
rect 3234 1264 3238 1301
rect 3254 1299 3261 1336
rect 3295 1313 3299 1356
rect 3315 1314 3319 1396
rect 3329 1337 3333 1396
rect 3349 1356 3353 1396
rect 3361 1390 3365 1396
rect 3355 1344 3358 1356
rect 3329 1329 3338 1337
rect 3254 1274 3261 1287
rect 3242 1268 3261 1274
rect 3242 1264 3246 1268
rect 3295 1264 3299 1301
rect 3315 1244 3319 1302
rect 3334 1300 3338 1329
rect 3354 1280 3358 1344
rect 3325 1276 3358 1280
rect 3325 1244 3329 1276
rect 3363 1268 3367 1378
rect 3381 1370 3385 1396
rect 3427 1392 3431 1396
rect 3395 1390 3431 1392
rect 3407 1388 3431 1390
rect 3349 1256 3351 1268
rect 3347 1244 3351 1256
rect 3357 1256 3359 1268
rect 3357 1244 3361 1256
rect 3379 1244 3383 1358
rect 3395 1252 3399 1378
rect 3435 1364 3439 1396
rect 3455 1376 3459 1416
rect 3463 1393 3467 1416
rect 3463 1386 3471 1393
rect 3433 1269 3439 1364
rect 3467 1357 3471 1386
rect 3463 1351 3471 1357
rect 3463 1305 3467 1351
rect 3485 1344 3489 1356
rect 3487 1332 3489 1344
rect 3433 1265 3457 1269
rect 3419 1260 3437 1261
rect 3407 1256 3437 1260
rect 3395 1248 3429 1252
rect 3425 1244 3429 1248
rect 3433 1244 3437 1256
rect 3453 1244 3457 1265
rect 3463 1244 3467 1293
rect 3485 1264 3489 1332
rect 3545 1313 3549 1396
rect 3617 1333 3621 1356
rect 3606 1321 3621 1333
rect 3625 1333 3629 1356
rect 3697 1333 3701 1356
rect 3625 1321 3634 1333
rect 3686 1321 3701 1333
rect 3705 1333 3709 1356
rect 3705 1321 3714 1333
rect 3545 1301 3554 1313
rect 3545 1244 3549 1301
rect 3605 1244 3609 1321
rect 3625 1244 3629 1321
rect 3685 1244 3689 1321
rect 3705 1244 3709 1321
rect 3751 1313 3755 1396
rect 3833 1393 3837 1416
rect 3829 1386 3837 1393
rect 3829 1357 3833 1386
rect 3841 1376 3845 1416
rect 3861 1364 3865 1396
rect 3869 1392 3873 1396
rect 3869 1390 3905 1392
rect 3869 1388 3893 1390
rect 3746 1301 3755 1313
rect 3751 1244 3755 1301
rect 3811 1344 3815 1356
rect 3829 1351 3837 1357
rect 3811 1332 3813 1344
rect 3811 1264 3815 1332
rect 3833 1305 3837 1351
rect 3833 1244 3837 1293
rect 3861 1269 3867 1364
rect 3843 1265 3867 1269
rect 3843 1244 3847 1265
rect 3863 1260 3881 1261
rect 3863 1256 3893 1260
rect 3863 1244 3867 1256
rect 3901 1252 3905 1378
rect 3915 1370 3919 1396
rect 3935 1390 3939 1396
rect 3871 1248 3905 1252
rect 3871 1244 3875 1248
rect 3917 1244 3921 1358
rect 3933 1268 3937 1378
rect 3947 1356 3951 1396
rect 3942 1344 3945 1356
rect 3942 1280 3946 1344
rect 3967 1337 3971 1396
rect 3962 1329 3971 1337
rect 3962 1300 3966 1329
rect 3981 1314 3985 1396
rect 4001 1313 4005 1356
rect 4056 1352 4060 1356
rect 4042 1344 4060 1352
rect 4042 1333 4046 1344
rect 3942 1276 3975 1280
rect 3941 1256 3943 1268
rect 3939 1244 3943 1256
rect 3949 1256 3951 1268
rect 3949 1244 3953 1256
rect 3971 1244 3975 1276
rect 3981 1244 3985 1302
rect 4001 1264 4005 1301
rect 4042 1276 4046 1321
rect 4064 1299 4068 1356
rect 4086 1353 4090 1396
rect 4086 1341 4093 1353
rect 4066 1287 4075 1299
rect 4042 1269 4055 1276
rect 4051 1264 4055 1269
rect 4071 1264 4075 1287
rect 4091 1264 4095 1341
rect 4151 1319 4155 1396
rect 4146 1307 4155 1319
rect 4149 1291 4155 1307
rect 4171 1319 4175 1396
rect 4243 1350 4247 1356
rect 4243 1338 4245 1350
rect 4265 1333 4269 1396
rect 4265 1321 4274 1333
rect 4171 1307 4174 1319
rect 4171 1291 4177 1307
rect 4149 1284 4157 1291
rect 4153 1264 4157 1284
rect 4163 1284 4177 1291
rect 4163 1264 4167 1284
rect 4243 1270 4245 1282
rect 4243 1264 4247 1270
rect 4265 1244 4269 1321
rect 4325 1319 4329 1396
rect 4326 1307 4329 1319
rect 4323 1291 4329 1307
rect 4345 1319 4349 1396
rect 4410 1353 4414 1396
rect 4407 1341 4414 1353
rect 4345 1307 4354 1319
rect 4345 1291 4351 1307
rect 4323 1284 4337 1291
rect 4333 1264 4337 1284
rect 4343 1284 4351 1291
rect 4343 1264 4347 1284
rect 4405 1264 4409 1341
rect 4432 1299 4436 1356
rect 4440 1352 4444 1356
rect 4510 1353 4514 1396
rect 4440 1344 4458 1352
rect 4454 1333 4458 1344
rect 4507 1341 4514 1353
rect 4425 1287 4434 1299
rect 4425 1264 4429 1287
rect 4454 1276 4458 1321
rect 4445 1269 4458 1276
rect 4445 1264 4449 1269
rect 4505 1264 4509 1341
rect 4532 1299 4536 1356
rect 4540 1352 4544 1356
rect 4540 1344 4558 1352
rect 4554 1333 4558 1344
rect 4591 1333 4595 1356
rect 4586 1321 4595 1333
rect 4599 1333 4603 1356
rect 4599 1321 4614 1333
rect 4525 1287 4534 1299
rect 4525 1264 4529 1287
rect 4554 1276 4558 1321
rect 4545 1269 4558 1276
rect 4545 1264 4549 1269
rect 4591 1244 4595 1321
rect 4611 1244 4615 1321
rect 4671 1313 4675 1396
rect 4666 1301 4675 1313
rect 4671 1244 4675 1301
rect 4745 1313 4749 1396
rect 4745 1301 4754 1313
rect 4745 1244 4749 1301
rect 52 1220 56 1224
rect 74 1220 78 1224
rect 82 1220 86 1224
rect 132 1220 136 1224
rect 140 1220 144 1224
rect 148 1220 152 1224
rect 232 1220 236 1224
rect 240 1220 244 1224
rect 248 1220 252 1224
rect 353 1220 357 1224
rect 363 1220 367 1224
rect 411 1220 415 1224
rect 431 1220 435 1224
rect 451 1220 455 1224
rect 514 1220 518 1224
rect 522 1220 526 1224
rect 544 1220 548 1224
rect 611 1220 615 1224
rect 631 1220 635 1224
rect 651 1220 655 1224
rect 711 1220 715 1224
rect 731 1220 735 1224
rect 751 1220 755 1224
rect 811 1220 815 1224
rect 821 1220 825 1224
rect 841 1220 845 1224
rect 933 1220 937 1224
rect 943 1220 947 1224
rect 993 1220 997 1224
rect 1003 1220 1007 1224
rect 1108 1220 1112 1224
rect 1116 1220 1120 1224
rect 1124 1220 1128 1224
rect 1185 1220 1189 1224
rect 1255 1220 1259 1224
rect 1275 1220 1279 1224
rect 1285 1220 1289 1224
rect 1331 1220 1335 1224
rect 1351 1220 1355 1224
rect 1371 1220 1375 1224
rect 1445 1220 1449 1224
rect 1465 1220 1469 1224
rect 1485 1220 1489 1224
rect 1533 1220 1537 1224
rect 1543 1220 1547 1224
rect 1611 1220 1615 1224
rect 1631 1220 1635 1224
rect 1651 1220 1655 1224
rect 1713 1220 1717 1224
rect 1723 1220 1727 1224
rect 1794 1220 1798 1224
rect 1802 1220 1806 1224
rect 1824 1220 1828 1224
rect 1892 1220 1896 1224
rect 1900 1220 1904 1224
rect 1908 1220 1912 1224
rect 1991 1220 1995 1224
rect 2011 1220 2015 1224
rect 2031 1220 2035 1224
rect 2091 1220 2095 1224
rect 2152 1220 2156 1224
rect 2160 1220 2164 1224
rect 2168 1220 2172 1224
rect 2253 1220 2257 1224
rect 2263 1220 2267 1224
rect 2331 1220 2335 1224
rect 2351 1220 2355 1224
rect 2371 1220 2375 1224
rect 2453 1220 2457 1224
rect 2463 1220 2467 1224
rect 2511 1220 2515 1224
rect 2583 1220 2587 1224
rect 2605 1220 2609 1224
rect 2651 1220 2655 1224
rect 2671 1220 2675 1224
rect 2691 1220 2695 1224
rect 2765 1220 2769 1224
rect 2785 1220 2789 1224
rect 2805 1220 2809 1224
rect 2825 1220 2829 1224
rect 2875 1220 2879 1224
rect 2895 1220 2899 1224
rect 2905 1220 2909 1224
rect 2927 1220 2931 1224
rect 2937 1220 2941 1224
rect 2959 1220 2963 1224
rect 3005 1220 3009 1224
rect 3013 1220 3017 1224
rect 3033 1220 3037 1224
rect 3043 1220 3047 1224
rect 3065 1220 3069 1224
rect 3125 1220 3129 1224
rect 3145 1220 3149 1224
rect 3212 1220 3216 1224
rect 3234 1220 3238 1224
rect 3242 1220 3246 1224
rect 3295 1220 3299 1224
rect 3315 1220 3319 1224
rect 3325 1220 3329 1224
rect 3347 1220 3351 1224
rect 3357 1220 3361 1224
rect 3379 1220 3383 1224
rect 3425 1220 3429 1224
rect 3433 1220 3437 1224
rect 3453 1220 3457 1224
rect 3463 1220 3467 1224
rect 3485 1220 3489 1224
rect 3545 1220 3549 1224
rect 3605 1220 3609 1224
rect 3625 1220 3629 1224
rect 3685 1220 3689 1224
rect 3705 1220 3709 1224
rect 3751 1220 3755 1224
rect 3811 1220 3815 1224
rect 3833 1220 3837 1224
rect 3843 1220 3847 1224
rect 3863 1220 3867 1224
rect 3871 1220 3875 1224
rect 3917 1220 3921 1224
rect 3939 1220 3943 1224
rect 3949 1220 3953 1224
rect 3971 1220 3975 1224
rect 3981 1220 3985 1224
rect 4001 1220 4005 1224
rect 4051 1220 4055 1224
rect 4071 1220 4075 1224
rect 4091 1220 4095 1224
rect 4153 1220 4157 1224
rect 4163 1220 4167 1224
rect 4243 1220 4247 1224
rect 4265 1220 4269 1224
rect 4333 1220 4337 1224
rect 4343 1220 4347 1224
rect 4405 1220 4409 1224
rect 4425 1220 4429 1224
rect 4445 1220 4449 1224
rect 4505 1220 4509 1224
rect 4525 1220 4529 1224
rect 4545 1220 4549 1224
rect 4591 1220 4595 1224
rect 4611 1220 4615 1224
rect 4671 1220 4675 1224
rect 4745 1220 4749 1224
rect 45 1196 49 1200
rect 65 1196 69 1200
rect 85 1196 89 1200
rect 131 1196 135 1200
rect 151 1196 155 1200
rect 171 1196 175 1200
rect 232 1196 236 1200
rect 240 1196 244 1200
rect 248 1196 252 1200
rect 334 1196 338 1200
rect 342 1196 346 1200
rect 364 1196 368 1200
rect 432 1196 436 1200
rect 440 1196 444 1200
rect 448 1196 452 1200
rect 534 1196 538 1200
rect 542 1196 546 1200
rect 564 1196 568 1200
rect 653 1196 657 1200
rect 663 1196 667 1200
rect 735 1196 739 1200
rect 755 1196 759 1200
rect 765 1196 769 1200
rect 848 1196 852 1200
rect 856 1196 860 1200
rect 864 1196 868 1200
rect 925 1196 929 1200
rect 945 1196 949 1200
rect 965 1196 969 1200
rect 1011 1196 1015 1200
rect 1031 1196 1035 1200
rect 1051 1196 1055 1200
rect 1125 1196 1129 1200
rect 1145 1196 1149 1200
rect 1165 1196 1169 1200
rect 1233 1196 1237 1200
rect 1243 1196 1247 1200
rect 1315 1196 1319 1200
rect 1335 1196 1339 1200
rect 1345 1196 1349 1200
rect 1393 1196 1397 1200
rect 1403 1196 1407 1200
rect 1485 1196 1489 1200
rect 1553 1196 1557 1200
rect 1563 1196 1567 1200
rect 1633 1196 1637 1200
rect 1643 1196 1647 1200
rect 1692 1196 1696 1200
rect 1700 1196 1704 1200
rect 1708 1196 1712 1200
rect 1813 1196 1817 1200
rect 1823 1196 1827 1200
rect 1872 1196 1876 1200
rect 1880 1196 1884 1200
rect 1888 1196 1892 1200
rect 1973 1196 1977 1200
rect 1983 1196 1987 1200
rect 2086 1196 2090 1200
rect 2094 1196 2098 1200
rect 2114 1196 2118 1200
rect 2122 1196 2126 1200
rect 2208 1196 2212 1200
rect 2216 1196 2220 1200
rect 2224 1196 2228 1200
rect 2293 1196 2297 1200
rect 2303 1196 2307 1200
rect 2354 1196 2358 1200
rect 2362 1196 2366 1200
rect 2384 1196 2388 1200
rect 2465 1196 2469 1200
rect 2533 1196 2537 1200
rect 2543 1196 2547 1200
rect 2605 1196 2609 1200
rect 2625 1196 2629 1200
rect 2645 1196 2649 1200
rect 2665 1196 2669 1200
rect 2711 1196 2715 1200
rect 2733 1196 2737 1200
rect 2795 1196 2799 1200
rect 2815 1196 2819 1200
rect 2825 1196 2829 1200
rect 2847 1196 2851 1200
rect 2857 1196 2861 1200
rect 2879 1196 2883 1200
rect 2925 1196 2929 1200
rect 2933 1196 2937 1200
rect 2953 1196 2957 1200
rect 2963 1196 2967 1200
rect 2985 1196 2989 1200
rect 3033 1196 3037 1200
rect 3043 1196 3047 1200
rect 3125 1196 3129 1200
rect 3145 1196 3149 1200
rect 3165 1196 3169 1200
rect 3211 1196 3215 1200
rect 3231 1196 3235 1200
rect 3251 1196 3255 1200
rect 3271 1196 3275 1200
rect 3343 1196 3347 1200
rect 3365 1196 3369 1200
rect 3411 1196 3415 1200
rect 3433 1196 3437 1200
rect 3491 1196 3495 1200
rect 3511 1196 3515 1200
rect 3531 1196 3535 1200
rect 3551 1196 3555 1200
rect 3571 1196 3575 1200
rect 3591 1196 3595 1200
rect 3611 1196 3615 1200
rect 3631 1196 3635 1200
rect 3691 1196 3695 1200
rect 3711 1196 3715 1200
rect 3731 1196 3735 1200
rect 3751 1196 3755 1200
rect 3771 1196 3775 1200
rect 3791 1196 3795 1200
rect 3811 1196 3815 1200
rect 3831 1196 3835 1200
rect 3891 1196 3895 1200
rect 3913 1196 3917 1200
rect 3973 1196 3977 1200
rect 3983 1196 3987 1200
rect 4051 1196 4055 1200
rect 4073 1196 4077 1200
rect 4083 1196 4087 1200
rect 4103 1196 4107 1200
rect 4111 1196 4115 1200
rect 4157 1196 4161 1200
rect 4179 1196 4183 1200
rect 4189 1196 4193 1200
rect 4211 1196 4215 1200
rect 4221 1196 4225 1200
rect 4241 1196 4245 1200
rect 4293 1196 4297 1200
rect 4303 1196 4307 1200
rect 4371 1196 4375 1200
rect 4391 1196 4395 1200
rect 4411 1196 4415 1200
rect 4493 1196 4497 1200
rect 4503 1196 4507 1200
rect 4551 1196 4555 1200
rect 4571 1196 4575 1200
rect 4591 1196 4595 1200
rect 4652 1196 4656 1200
rect 4660 1196 4664 1200
rect 4668 1196 4672 1200
rect 45 1079 49 1156
rect 65 1133 69 1156
rect 85 1151 89 1156
rect 131 1151 135 1156
rect 85 1144 98 1151
rect 65 1121 74 1133
rect 47 1067 54 1079
rect 50 1024 54 1067
rect 72 1064 76 1121
rect 94 1099 98 1144
rect 122 1144 135 1151
rect 122 1099 126 1144
rect 151 1133 155 1156
rect 146 1121 155 1133
rect 94 1076 98 1087
rect 80 1068 98 1076
rect 122 1076 126 1087
rect 122 1068 140 1076
rect 80 1064 84 1068
rect 136 1064 140 1068
rect 144 1064 148 1121
rect 171 1079 175 1156
rect 334 1152 338 1156
rect 319 1146 338 1152
rect 232 1079 236 1136
rect 166 1067 173 1079
rect 226 1067 236 1079
rect 166 1024 170 1067
rect 220 1036 226 1067
rect 240 1059 244 1136
rect 248 1079 252 1136
rect 319 1133 326 1146
rect 319 1084 326 1121
rect 342 1119 346 1156
rect 364 1133 368 1176
rect 534 1152 538 1156
rect 519 1146 538 1152
rect 366 1121 375 1133
rect 340 1084 346 1107
rect 248 1067 255 1079
rect 267 1067 275 1079
rect 319 1078 335 1084
rect 340 1078 355 1084
rect 240 1040 246 1047
rect 240 1036 255 1040
rect 220 1032 235 1036
rect 231 1024 235 1032
rect 251 1024 255 1036
rect 271 1024 275 1067
rect 331 1064 335 1078
rect 351 1064 355 1078
rect 371 1064 375 1121
rect 432 1079 436 1136
rect 426 1067 436 1079
rect 420 1036 426 1067
rect 440 1059 444 1136
rect 448 1079 452 1136
rect 519 1133 526 1146
rect 519 1084 526 1121
rect 542 1119 546 1156
rect 564 1133 568 1176
rect 653 1136 657 1156
rect 566 1121 575 1133
rect 540 1084 546 1107
rect 448 1067 455 1079
rect 467 1067 475 1079
rect 519 1078 535 1084
rect 540 1078 555 1084
rect 440 1040 446 1047
rect 440 1036 455 1040
rect 420 1032 435 1036
rect 431 1024 435 1032
rect 451 1024 455 1036
rect 471 1024 475 1067
rect 531 1064 535 1078
rect 551 1064 555 1078
rect 571 1064 575 1121
rect 643 1129 657 1136
rect 663 1136 667 1156
rect 735 1150 739 1156
rect 721 1138 733 1150
rect 663 1129 671 1136
rect 643 1113 649 1129
rect 646 1101 649 1113
rect 645 1024 649 1101
rect 665 1113 671 1129
rect 665 1101 674 1113
rect 665 1024 669 1101
rect 721 1064 725 1138
rect 755 1113 759 1156
rect 746 1101 759 1113
rect 743 1024 747 1101
rect 765 1099 769 1156
rect 765 1087 774 1099
rect 765 1024 769 1087
rect 848 1079 852 1136
rect 825 1067 833 1079
rect 845 1067 852 1079
rect 825 1024 829 1067
rect 856 1059 860 1136
rect 864 1079 868 1136
rect 925 1079 929 1156
rect 945 1133 949 1156
rect 965 1151 969 1156
rect 1011 1151 1015 1156
rect 965 1144 978 1151
rect 945 1121 954 1133
rect 864 1067 874 1079
rect 927 1067 934 1079
rect 854 1040 860 1047
rect 845 1036 860 1040
rect 874 1036 880 1067
rect 845 1024 849 1036
rect 865 1032 880 1036
rect 865 1024 869 1032
rect 930 1024 934 1067
rect 952 1064 956 1121
rect 974 1099 978 1144
rect 1002 1144 1015 1151
rect 1002 1099 1006 1144
rect 1031 1133 1035 1156
rect 1026 1121 1035 1133
rect 974 1076 978 1087
rect 960 1068 978 1076
rect 1002 1076 1006 1087
rect 1002 1068 1020 1076
rect 960 1064 964 1068
rect 1016 1064 1020 1068
rect 1024 1064 1028 1121
rect 1051 1079 1055 1156
rect 1125 1079 1129 1156
rect 1145 1133 1149 1156
rect 1165 1151 1169 1156
rect 1165 1144 1178 1151
rect 1145 1121 1154 1133
rect 1046 1067 1053 1079
rect 1127 1067 1134 1079
rect 1046 1024 1050 1067
rect 1130 1024 1134 1067
rect 1152 1064 1156 1121
rect 1174 1099 1178 1144
rect 1233 1136 1237 1156
rect 1223 1129 1237 1136
rect 1243 1136 1247 1156
rect 1315 1150 1319 1156
rect 1301 1138 1313 1150
rect 1243 1129 1251 1136
rect 1223 1113 1229 1129
rect 1226 1101 1229 1113
rect 1174 1076 1178 1087
rect 1160 1068 1178 1076
rect 1160 1064 1164 1068
rect 1225 1024 1229 1101
rect 1245 1113 1251 1129
rect 1245 1101 1254 1113
rect 1245 1024 1249 1101
rect 1301 1064 1305 1138
rect 1335 1113 1339 1156
rect 1326 1101 1339 1113
rect 1323 1024 1327 1101
rect 1345 1099 1349 1156
rect 1393 1136 1397 1156
rect 1389 1129 1397 1136
rect 1403 1136 1407 1156
rect 1403 1129 1417 1136
rect 1389 1113 1395 1129
rect 1386 1101 1395 1113
rect 1345 1087 1354 1099
rect 1345 1024 1349 1087
rect 1391 1024 1395 1101
rect 1411 1113 1417 1129
rect 1485 1133 1489 1156
rect 1553 1136 1557 1156
rect 1485 1121 1494 1133
rect 1543 1129 1557 1136
rect 1563 1136 1567 1156
rect 1633 1136 1637 1156
rect 1563 1129 1571 1136
rect 1411 1101 1414 1113
rect 1411 1024 1415 1101
rect 1485 1064 1489 1121
rect 1543 1113 1549 1129
rect 1546 1101 1549 1113
rect 1545 1024 1549 1101
rect 1565 1113 1571 1129
rect 1623 1129 1637 1136
rect 1643 1136 1647 1156
rect 1813 1136 1817 1156
rect 1643 1129 1651 1136
rect 1623 1113 1629 1129
rect 1565 1101 1574 1113
rect 1626 1101 1629 1113
rect 1565 1024 1569 1101
rect 1625 1024 1629 1101
rect 1645 1113 1651 1129
rect 1645 1101 1654 1113
rect 1645 1024 1649 1101
rect 1692 1079 1696 1136
rect 1686 1067 1696 1079
rect 1680 1036 1686 1067
rect 1700 1059 1704 1136
rect 1708 1079 1712 1136
rect 1803 1129 1817 1136
rect 1823 1136 1827 1156
rect 1973 1136 1977 1156
rect 1823 1129 1831 1136
rect 1803 1113 1809 1129
rect 1806 1101 1809 1113
rect 1708 1067 1715 1079
rect 1727 1067 1735 1079
rect 1700 1040 1706 1047
rect 1700 1036 1715 1040
rect 1680 1032 1695 1036
rect 1691 1024 1695 1032
rect 1711 1024 1715 1036
rect 1731 1024 1735 1067
rect 1805 1024 1809 1101
rect 1825 1113 1831 1129
rect 1825 1101 1834 1113
rect 1825 1024 1829 1101
rect 1872 1079 1876 1136
rect 1866 1067 1876 1079
rect 1860 1036 1866 1067
rect 1880 1059 1884 1136
rect 1888 1079 1892 1136
rect 1969 1129 1977 1136
rect 1983 1136 1987 1156
rect 2086 1151 2090 1156
rect 2060 1147 2090 1151
rect 1983 1129 1997 1136
rect 1969 1113 1975 1129
rect 1966 1101 1975 1113
rect 1888 1067 1895 1079
rect 1907 1067 1915 1079
rect 1880 1040 1886 1047
rect 1880 1036 1895 1040
rect 1860 1032 1875 1036
rect 1871 1024 1875 1032
rect 1891 1024 1895 1036
rect 1911 1024 1915 1067
rect 1971 1024 1975 1101
rect 1991 1113 1997 1129
rect 1991 1101 1994 1113
rect 1991 1024 1995 1101
rect 2060 1099 2066 1147
rect 2094 1142 2098 1156
rect 2085 1135 2098 1142
rect 2085 1133 2089 1135
rect 2114 1133 2118 1156
rect 2122 1148 2126 1156
rect 2122 1141 2139 1148
rect 2087 1121 2089 1133
rect 2066 1087 2069 1099
rect 2065 1064 2069 1087
rect 2085 1064 2089 1121
rect 2114 1092 2118 1121
rect 2133 1099 2139 1141
rect 2293 1136 2297 1156
rect 2105 1086 2118 1092
rect 2125 1087 2133 1092
rect 2125 1086 2145 1087
rect 2105 1064 2109 1086
rect 2125 1064 2129 1086
rect 2208 1079 2212 1136
rect 2185 1067 2193 1079
rect 2205 1067 2212 1079
rect 2185 1024 2189 1067
rect 2216 1059 2220 1136
rect 2224 1079 2228 1136
rect 2283 1129 2297 1136
rect 2303 1136 2307 1156
rect 2354 1152 2358 1156
rect 2339 1146 2358 1152
rect 2303 1129 2311 1136
rect 2339 1133 2346 1146
rect 2283 1113 2289 1129
rect 2286 1101 2289 1113
rect 2224 1067 2234 1079
rect 2214 1040 2220 1047
rect 2205 1036 2220 1040
rect 2234 1036 2240 1067
rect 2205 1024 2209 1036
rect 2225 1032 2240 1036
rect 2225 1024 2229 1032
rect 2285 1024 2289 1101
rect 2305 1113 2311 1129
rect 2305 1101 2314 1113
rect 2305 1024 2309 1101
rect 2339 1084 2346 1121
rect 2362 1119 2366 1156
rect 2384 1133 2388 1176
rect 2386 1121 2395 1133
rect 2360 1084 2366 1107
rect 2339 1078 2355 1084
rect 2360 1078 2375 1084
rect 2351 1064 2355 1078
rect 2371 1064 2375 1078
rect 2391 1064 2395 1121
rect 2465 1119 2469 1176
rect 2533 1136 2537 1156
rect 2523 1129 2537 1136
rect 2543 1136 2547 1156
rect 2543 1129 2551 1136
rect 2465 1107 2474 1119
rect 2523 1113 2529 1129
rect 2465 1024 2469 1107
rect 2526 1101 2529 1113
rect 2525 1024 2529 1101
rect 2545 1113 2551 1129
rect 2545 1101 2554 1113
rect 2545 1024 2549 1101
rect 2605 1099 2609 1156
rect 2625 1133 2629 1156
rect 2645 1133 2649 1156
rect 2665 1149 2669 1156
rect 2665 1145 2680 1149
rect 2645 1121 2654 1133
rect 2607 1087 2609 1099
rect 2605 1072 2609 1087
rect 2605 1068 2619 1072
rect 2615 1064 2619 1068
rect 2625 1064 2629 1121
rect 2645 1072 2651 1121
rect 2674 1099 2680 1145
rect 2711 1099 2715 1176
rect 2733 1150 2737 1156
rect 2735 1138 2737 1150
rect 2795 1119 2799 1156
rect 2815 1118 2819 1176
rect 2825 1144 2829 1176
rect 2847 1164 2851 1176
rect 2849 1152 2851 1164
rect 2857 1164 2861 1176
rect 2857 1152 2859 1164
rect 2825 1140 2858 1144
rect 2706 1087 2715 1099
rect 2674 1072 2679 1087
rect 2645 1068 2659 1072
rect 2655 1064 2659 1068
rect 2665 1068 2679 1072
rect 2665 1064 2669 1068
rect 2711 1024 2715 1087
rect 2735 1070 2737 1082
rect 2733 1064 2737 1070
rect 2795 1064 2799 1107
rect 2815 1024 2819 1106
rect 2834 1091 2838 1120
rect 2829 1083 2838 1091
rect 2829 1024 2833 1083
rect 2854 1076 2858 1140
rect 2855 1064 2858 1076
rect 2849 1024 2853 1064
rect 2863 1042 2867 1152
rect 2879 1062 2883 1176
rect 2925 1172 2929 1176
rect 2895 1168 2929 1172
rect 2861 1024 2865 1030
rect 2881 1024 2885 1050
rect 2895 1042 2899 1168
rect 2933 1164 2937 1176
rect 2907 1160 2937 1164
rect 2919 1159 2937 1160
rect 2953 1155 2957 1176
rect 2933 1151 2957 1155
rect 2933 1056 2939 1151
rect 2963 1127 2967 1176
rect 2963 1069 2967 1115
rect 2985 1088 2989 1156
rect 3033 1136 3037 1156
rect 3029 1129 3037 1136
rect 3043 1136 3047 1156
rect 3043 1129 3057 1136
rect 3029 1113 3035 1129
rect 3026 1101 3035 1113
rect 2987 1076 2989 1088
rect 2963 1063 2971 1069
rect 2985 1064 2989 1076
rect 2907 1030 2931 1032
rect 2895 1028 2931 1030
rect 2927 1024 2931 1028
rect 2935 1024 2939 1056
rect 2955 1004 2959 1044
rect 2967 1034 2971 1063
rect 2963 1027 2971 1034
rect 2963 1004 2967 1027
rect 3031 1024 3035 1101
rect 3051 1113 3057 1129
rect 3051 1101 3054 1113
rect 3051 1024 3055 1101
rect 3125 1079 3129 1156
rect 3145 1133 3149 1156
rect 3165 1151 3169 1156
rect 3211 1152 3215 1156
rect 3231 1152 3235 1156
rect 3251 1152 3255 1156
rect 3271 1152 3275 1156
rect 3165 1144 3178 1151
rect 3145 1121 3154 1133
rect 3127 1067 3134 1079
rect 3130 1024 3134 1067
rect 3152 1064 3156 1121
rect 3174 1099 3178 1144
rect 3211 1148 3275 1152
rect 3343 1150 3347 1156
rect 3211 1099 3217 1148
rect 3343 1138 3345 1150
rect 3365 1099 3369 1176
rect 3411 1099 3415 1176
rect 3433 1150 3437 1156
rect 3435 1138 3437 1150
rect 3211 1087 3214 1099
rect 3365 1087 3374 1099
rect 3406 1087 3415 1099
rect 3174 1076 3178 1087
rect 3160 1068 3178 1076
rect 3211 1072 3217 1087
rect 3211 1068 3275 1072
rect 3160 1064 3164 1068
rect 3211 1064 3215 1068
rect 3231 1064 3235 1068
rect 3251 1064 3255 1068
rect 3271 1064 3275 1068
rect 3343 1070 3345 1082
rect 3343 1064 3347 1070
rect 3365 1024 3369 1087
rect 3411 1024 3415 1087
rect 3491 1133 3495 1156
rect 3511 1133 3515 1156
rect 3531 1136 3535 1156
rect 3551 1136 3555 1156
rect 3571 1136 3575 1156
rect 3591 1136 3595 1156
rect 3611 1136 3615 1156
rect 3631 1136 3635 1156
rect 3491 1121 3494 1133
rect 3506 1121 3515 1133
rect 3542 1124 3555 1136
rect 3582 1124 3595 1136
rect 3622 1124 3635 1136
rect 3435 1070 3437 1082
rect 3433 1064 3437 1070
rect 3491 1064 3495 1121
rect 3511 1064 3515 1121
rect 3531 1064 3535 1124
rect 3551 1064 3555 1124
rect 3571 1064 3575 1124
rect 3591 1064 3595 1124
rect 3611 1064 3615 1124
rect 3631 1064 3635 1124
rect 3691 1133 3695 1156
rect 3711 1133 3715 1156
rect 3731 1136 3735 1156
rect 3751 1136 3755 1156
rect 3771 1136 3775 1156
rect 3791 1136 3795 1156
rect 3811 1136 3815 1156
rect 3831 1136 3835 1156
rect 3691 1121 3694 1133
rect 3706 1121 3715 1133
rect 3742 1124 3755 1136
rect 3782 1124 3795 1136
rect 3822 1124 3835 1136
rect 3691 1064 3695 1121
rect 3711 1064 3715 1121
rect 3731 1064 3735 1124
rect 3751 1064 3755 1124
rect 3771 1064 3775 1124
rect 3791 1064 3795 1124
rect 3811 1064 3815 1124
rect 3831 1064 3835 1124
rect 3891 1099 3895 1176
rect 3913 1150 3917 1156
rect 3915 1138 3917 1150
rect 3973 1136 3977 1156
rect 3969 1129 3977 1136
rect 3983 1136 3987 1156
rect 3983 1129 3997 1136
rect 3969 1113 3975 1129
rect 3966 1101 3975 1113
rect 3886 1087 3895 1099
rect 3891 1024 3895 1087
rect 3915 1070 3917 1082
rect 3913 1064 3917 1070
rect 3971 1024 3975 1101
rect 3991 1113 3997 1129
rect 3991 1101 3994 1113
rect 3991 1024 3995 1101
rect 4051 1088 4055 1156
rect 4073 1127 4077 1176
rect 4083 1155 4087 1176
rect 4103 1164 4107 1176
rect 4111 1172 4115 1176
rect 4111 1168 4145 1172
rect 4103 1160 4133 1164
rect 4103 1159 4121 1160
rect 4083 1151 4107 1155
rect 4051 1076 4053 1088
rect 4051 1064 4055 1076
rect 4073 1069 4077 1115
rect 4069 1063 4077 1069
rect 4069 1034 4073 1063
rect 4101 1056 4107 1151
rect 4069 1027 4077 1034
rect 4073 1004 4077 1027
rect 4081 1004 4085 1044
rect 4101 1024 4105 1056
rect 4141 1042 4145 1168
rect 4157 1062 4161 1176
rect 4179 1164 4183 1176
rect 4181 1152 4183 1164
rect 4189 1164 4193 1176
rect 4189 1152 4191 1164
rect 4109 1030 4133 1032
rect 4109 1028 4145 1030
rect 4109 1024 4113 1028
rect 4155 1024 4159 1050
rect 4173 1042 4177 1152
rect 4211 1144 4215 1176
rect 4182 1140 4215 1144
rect 4182 1076 4186 1140
rect 4202 1091 4206 1120
rect 4221 1118 4225 1176
rect 4241 1119 4245 1156
rect 4293 1136 4297 1156
rect 4289 1129 4297 1136
rect 4303 1136 4307 1156
rect 4371 1151 4375 1156
rect 4362 1144 4375 1151
rect 4303 1129 4317 1136
rect 4289 1113 4295 1129
rect 4202 1083 4211 1091
rect 4182 1064 4185 1076
rect 4175 1024 4179 1030
rect 4187 1024 4191 1064
rect 4207 1024 4211 1083
rect 4221 1024 4225 1106
rect 4241 1064 4245 1107
rect 4286 1101 4295 1113
rect 4291 1024 4295 1101
rect 4311 1113 4317 1129
rect 4311 1101 4314 1113
rect 4311 1024 4315 1101
rect 4362 1099 4366 1144
rect 4391 1133 4395 1156
rect 4386 1121 4395 1133
rect 4362 1076 4366 1087
rect 4362 1068 4380 1076
rect 4376 1064 4380 1068
rect 4384 1064 4388 1121
rect 4411 1079 4415 1156
rect 4493 1136 4497 1156
rect 4483 1129 4497 1136
rect 4503 1136 4507 1156
rect 4551 1151 4555 1156
rect 4542 1144 4555 1151
rect 4503 1129 4511 1136
rect 4483 1113 4489 1129
rect 4486 1101 4489 1113
rect 4406 1067 4413 1079
rect 4406 1024 4410 1067
rect 4485 1024 4489 1101
rect 4505 1113 4511 1129
rect 4505 1101 4514 1113
rect 4505 1024 4509 1101
rect 4542 1099 4546 1144
rect 4571 1133 4575 1156
rect 4566 1121 4575 1133
rect 4542 1076 4546 1087
rect 4542 1068 4560 1076
rect 4556 1064 4560 1068
rect 4564 1064 4568 1121
rect 4591 1079 4595 1156
rect 4652 1079 4656 1136
rect 4586 1067 4593 1079
rect 4646 1067 4656 1079
rect 4586 1024 4590 1067
rect 4640 1036 4646 1067
rect 4660 1059 4664 1136
rect 4668 1079 4672 1136
rect 4668 1067 4675 1079
rect 4687 1067 4695 1079
rect 4660 1040 4666 1047
rect 4660 1036 4675 1040
rect 4640 1032 4655 1036
rect 4651 1024 4655 1032
rect 4671 1024 4675 1036
rect 4691 1024 4695 1067
rect 50 980 54 984
rect 72 980 76 984
rect 80 980 84 984
rect 136 980 140 984
rect 144 980 148 984
rect 166 980 170 984
rect 231 980 235 984
rect 251 980 255 984
rect 271 980 275 984
rect 331 980 335 984
rect 351 980 355 984
rect 371 980 375 984
rect 431 980 435 984
rect 451 980 455 984
rect 471 980 475 984
rect 531 980 535 984
rect 551 980 555 984
rect 571 980 575 984
rect 645 980 649 984
rect 665 980 669 984
rect 721 980 725 984
rect 743 980 747 984
rect 765 980 769 984
rect 825 980 829 984
rect 845 980 849 984
rect 865 980 869 984
rect 930 980 934 984
rect 952 980 956 984
rect 960 980 964 984
rect 1016 980 1020 984
rect 1024 980 1028 984
rect 1046 980 1050 984
rect 1130 980 1134 984
rect 1152 980 1156 984
rect 1160 980 1164 984
rect 1225 980 1229 984
rect 1245 980 1249 984
rect 1301 980 1305 984
rect 1323 980 1327 984
rect 1345 980 1349 984
rect 1391 980 1395 984
rect 1411 980 1415 984
rect 1485 980 1489 984
rect 1545 980 1549 984
rect 1565 980 1569 984
rect 1625 980 1629 984
rect 1645 980 1649 984
rect 1691 980 1695 984
rect 1711 980 1715 984
rect 1731 980 1735 984
rect 1805 980 1809 984
rect 1825 980 1829 984
rect 1871 980 1875 984
rect 1891 980 1895 984
rect 1911 980 1915 984
rect 1971 980 1975 984
rect 1991 980 1995 984
rect 2065 980 2069 984
rect 2085 980 2089 984
rect 2105 980 2109 984
rect 2125 980 2129 984
rect 2185 980 2189 984
rect 2205 980 2209 984
rect 2225 980 2229 984
rect 2285 980 2289 984
rect 2305 980 2309 984
rect 2351 980 2355 984
rect 2371 980 2375 984
rect 2391 980 2395 984
rect 2465 980 2469 984
rect 2525 980 2529 984
rect 2545 980 2549 984
rect 2615 980 2619 984
rect 2625 980 2629 984
rect 2655 980 2659 984
rect 2665 980 2669 984
rect 2711 980 2715 984
rect 2733 980 2737 984
rect 2795 980 2799 984
rect 2815 980 2819 984
rect 2829 980 2833 984
rect 2849 980 2853 984
rect 2861 980 2865 984
rect 2881 980 2885 984
rect 2927 980 2931 984
rect 2935 980 2939 984
rect 2955 980 2959 984
rect 2963 980 2967 984
rect 2985 980 2989 984
rect 3031 980 3035 984
rect 3051 980 3055 984
rect 3130 980 3134 984
rect 3152 980 3156 984
rect 3160 980 3164 984
rect 3211 980 3215 984
rect 3231 980 3235 984
rect 3251 980 3255 984
rect 3271 980 3275 984
rect 3343 980 3347 984
rect 3365 980 3369 984
rect 3411 980 3415 984
rect 3433 980 3437 984
rect 3491 980 3495 984
rect 3511 980 3515 984
rect 3531 980 3535 984
rect 3551 980 3555 984
rect 3571 980 3575 984
rect 3591 980 3595 984
rect 3611 980 3615 984
rect 3631 980 3635 984
rect 3691 980 3695 984
rect 3711 980 3715 984
rect 3731 980 3735 984
rect 3751 980 3755 984
rect 3771 980 3775 984
rect 3791 980 3795 984
rect 3811 980 3815 984
rect 3831 980 3835 984
rect 3891 980 3895 984
rect 3913 980 3917 984
rect 3971 980 3975 984
rect 3991 980 3995 984
rect 4051 980 4055 984
rect 4073 980 4077 984
rect 4081 980 4085 984
rect 4101 980 4105 984
rect 4109 980 4113 984
rect 4155 980 4159 984
rect 4175 980 4179 984
rect 4187 980 4191 984
rect 4207 980 4211 984
rect 4221 980 4225 984
rect 4241 980 4245 984
rect 4291 980 4295 984
rect 4311 980 4315 984
rect 4376 980 4380 984
rect 4384 980 4388 984
rect 4406 980 4410 984
rect 4485 980 4489 984
rect 4505 980 4509 984
rect 4556 980 4560 984
rect 4564 980 4568 984
rect 4586 980 4590 984
rect 4651 980 4655 984
rect 4671 980 4675 984
rect 4691 980 4695 984
rect 45 956 49 960
rect 65 956 69 960
rect 121 956 125 960
rect 143 956 147 960
rect 165 956 169 960
rect 230 956 234 960
rect 252 956 256 960
rect 260 956 264 960
rect 325 956 329 960
rect 345 956 349 960
rect 365 956 369 960
rect 385 956 389 960
rect 443 956 447 960
rect 465 956 469 960
rect 511 956 515 960
rect 585 956 589 960
rect 645 956 649 960
rect 665 956 669 960
rect 685 956 689 960
rect 731 956 735 960
rect 751 956 755 960
rect 771 956 775 960
rect 841 956 845 960
rect 863 956 867 960
rect 885 956 889 960
rect 931 956 935 960
rect 951 956 955 960
rect 1025 956 1029 960
rect 1045 956 1049 960
rect 1065 956 1069 960
rect 1116 956 1120 960
rect 1124 956 1128 960
rect 1146 956 1150 960
rect 1225 956 1229 960
rect 1245 956 1249 960
rect 1265 956 1269 960
rect 1311 956 1315 960
rect 1376 956 1380 960
rect 1384 956 1388 960
rect 1406 956 1410 960
rect 1485 956 1489 960
rect 1505 956 1509 960
rect 1551 956 1555 960
rect 1571 956 1575 960
rect 1650 956 1654 960
rect 1672 956 1676 960
rect 1680 956 1684 960
rect 1731 956 1735 960
rect 1753 956 1757 960
rect 1775 956 1779 960
rect 1845 956 1849 960
rect 1905 956 1909 960
rect 1925 956 1929 960
rect 1971 956 1975 960
rect 2045 956 2049 960
rect 2065 956 2069 960
rect 2085 956 2089 960
rect 2131 956 2135 960
rect 2196 956 2200 960
rect 2204 956 2208 960
rect 2226 956 2230 960
rect 2305 956 2309 960
rect 2325 956 2329 960
rect 2345 956 2349 960
rect 2391 956 2395 960
rect 2451 956 2455 960
rect 2471 956 2475 960
rect 2491 956 2495 960
rect 2565 956 2569 960
rect 2585 956 2589 960
rect 2605 956 2609 960
rect 2651 956 2655 960
rect 2671 956 2675 960
rect 2691 956 2695 960
rect 2765 956 2769 960
rect 2785 956 2789 960
rect 2855 956 2859 960
rect 2865 956 2869 960
rect 2895 956 2899 960
rect 2905 956 2909 960
rect 2965 956 2969 960
rect 3037 956 3041 960
rect 3045 956 3049 960
rect 3117 956 3121 960
rect 3125 956 3129 960
rect 3171 956 3175 960
rect 3236 956 3240 960
rect 3244 956 3248 960
rect 3266 956 3270 960
rect 3331 956 3335 960
rect 3351 956 3355 960
rect 3411 956 3415 960
rect 3433 956 3437 960
rect 3441 956 3445 960
rect 3461 956 3465 960
rect 3469 956 3473 960
rect 3515 956 3519 960
rect 3535 956 3539 960
rect 3547 956 3551 960
rect 3567 956 3571 960
rect 3581 956 3585 960
rect 3601 956 3605 960
rect 3651 956 3655 960
rect 3673 956 3677 960
rect 3735 956 3739 960
rect 3755 956 3759 960
rect 3769 956 3773 960
rect 3789 956 3793 960
rect 3801 956 3805 960
rect 3821 956 3825 960
rect 3867 956 3871 960
rect 3875 956 3879 960
rect 3895 956 3899 960
rect 3903 956 3907 960
rect 3925 956 3929 960
rect 3990 956 3994 960
rect 4012 956 4016 960
rect 4020 956 4024 960
rect 4071 956 4075 960
rect 4093 956 4097 960
rect 4101 956 4105 960
rect 4121 956 4125 960
rect 4129 956 4133 960
rect 4175 956 4179 960
rect 4195 956 4199 960
rect 4207 956 4211 960
rect 4227 956 4231 960
rect 4241 956 4245 960
rect 4261 956 4265 960
rect 4315 956 4319 960
rect 4335 956 4339 960
rect 4349 956 4353 960
rect 4369 956 4373 960
rect 4381 956 4385 960
rect 4401 956 4405 960
rect 4447 956 4451 960
rect 4455 956 4459 960
rect 4475 956 4479 960
rect 4483 956 4487 960
rect 4505 956 4509 960
rect 4556 956 4560 960
rect 4564 956 4568 960
rect 4586 956 4590 960
rect 4656 956 4660 960
rect 4664 956 4668 960
rect 4686 956 4690 960
rect 45 839 49 916
rect 46 827 49 839
rect 43 811 49 827
rect 65 839 69 916
rect 65 827 74 839
rect 65 811 71 827
rect 43 804 57 811
rect 53 784 57 804
rect 63 804 71 811
rect 63 784 67 804
rect 121 802 125 876
rect 143 839 147 916
rect 165 853 169 916
rect 230 873 234 916
rect 227 861 234 873
rect 165 841 174 853
rect 146 827 159 839
rect 121 790 133 802
rect 135 784 139 790
rect 155 784 159 827
rect 165 784 169 841
rect 225 784 229 861
rect 252 819 256 876
rect 260 872 264 876
rect 260 864 278 872
rect 274 853 278 864
rect 325 853 329 876
rect 326 841 329 853
rect 245 807 254 819
rect 245 784 249 807
rect 274 796 278 841
rect 265 789 278 796
rect 320 793 326 841
rect 345 819 349 876
rect 365 854 369 876
rect 385 854 389 876
rect 443 870 447 876
rect 443 858 445 870
rect 365 848 378 854
rect 385 853 405 854
rect 385 848 393 853
rect 374 819 378 848
rect 465 853 469 916
rect 465 841 474 853
rect 347 807 349 819
rect 345 805 349 807
rect 345 798 358 805
rect 320 789 350 793
rect 265 784 269 789
rect 346 784 350 789
rect 354 784 358 798
rect 374 784 378 807
rect 393 799 399 841
rect 382 792 399 799
rect 382 784 386 792
rect 443 790 445 802
rect 443 784 447 790
rect 465 764 469 841
rect 511 833 515 916
rect 506 821 515 833
rect 511 764 515 821
rect 585 833 589 916
rect 731 908 735 916
rect 720 904 735 908
rect 751 904 755 916
rect 585 821 594 833
rect 585 764 589 821
rect 645 819 649 876
rect 665 862 669 876
rect 685 862 689 876
rect 720 873 726 904
rect 740 900 755 904
rect 740 893 746 900
rect 665 856 680 862
rect 685 856 701 862
rect 726 861 736 873
rect 674 833 680 856
rect 645 807 654 819
rect 652 764 656 807
rect 674 784 678 821
rect 694 819 701 856
rect 694 794 701 807
rect 732 804 736 861
rect 740 804 744 881
rect 771 873 775 916
rect 748 861 755 873
rect 767 861 775 873
rect 748 804 752 861
rect 682 788 701 794
rect 682 784 686 788
rect 841 802 845 876
rect 863 839 867 916
rect 885 853 889 916
rect 885 841 894 853
rect 866 827 879 839
rect 841 790 853 802
rect 855 784 859 790
rect 875 784 879 827
rect 885 784 889 841
rect 931 839 935 916
rect 926 827 935 839
rect 929 811 935 827
rect 951 839 955 916
rect 1025 873 1029 916
rect 1045 904 1049 916
rect 1065 908 1069 916
rect 1065 904 1080 908
rect 1045 900 1060 904
rect 1054 893 1060 900
rect 1025 861 1033 873
rect 1045 861 1052 873
rect 951 827 954 839
rect 951 811 957 827
rect 929 804 937 811
rect 933 784 937 804
rect 943 804 957 811
rect 1048 804 1052 861
rect 1056 804 1060 881
rect 1074 873 1080 904
rect 1064 861 1074 873
rect 1116 872 1120 876
rect 1102 864 1120 872
rect 1064 804 1068 861
rect 1102 853 1106 864
rect 943 784 947 804
rect 1102 796 1106 841
rect 1124 819 1128 876
rect 1146 873 1150 916
rect 1225 873 1229 916
rect 1245 904 1249 916
rect 1265 908 1269 916
rect 1265 904 1280 908
rect 1245 900 1260 904
rect 1254 893 1260 900
rect 1146 861 1153 873
rect 1225 861 1233 873
rect 1245 861 1252 873
rect 1126 807 1135 819
rect 1102 789 1115 796
rect 1111 784 1115 789
rect 1131 784 1135 807
rect 1151 784 1155 861
rect 1248 804 1252 861
rect 1256 804 1260 881
rect 1274 873 1280 904
rect 1264 861 1274 873
rect 1264 804 1268 861
rect 1311 833 1315 916
rect 1376 872 1380 876
rect 1362 864 1380 872
rect 1362 853 1366 864
rect 1306 821 1315 833
rect 1311 764 1315 821
rect 1362 796 1366 841
rect 1384 819 1388 876
rect 1406 873 1410 916
rect 1406 861 1413 873
rect 1386 807 1395 819
rect 1362 789 1375 796
rect 1371 784 1375 789
rect 1391 784 1395 807
rect 1411 784 1415 861
rect 1485 839 1489 916
rect 1486 827 1489 839
rect 1483 811 1489 827
rect 1505 839 1509 916
rect 1551 839 1555 916
rect 1505 827 1514 839
rect 1546 827 1555 839
rect 1505 811 1511 827
rect 1483 804 1497 811
rect 1493 784 1497 804
rect 1503 804 1511 811
rect 1549 811 1555 827
rect 1571 839 1575 916
rect 1650 873 1654 916
rect 1647 861 1654 873
rect 1571 827 1574 839
rect 1571 811 1577 827
rect 1549 804 1557 811
rect 1503 784 1507 804
rect 1553 784 1557 804
rect 1563 804 1577 811
rect 1563 784 1567 804
rect 1645 784 1649 861
rect 1672 819 1676 876
rect 1680 872 1684 876
rect 1680 864 1698 872
rect 1694 853 1698 864
rect 1731 853 1735 916
rect 1726 841 1735 853
rect 1665 807 1674 819
rect 1665 784 1669 807
rect 1694 796 1698 841
rect 1685 789 1698 796
rect 1685 784 1689 789
rect 1731 784 1735 841
rect 1753 839 1757 916
rect 1741 827 1754 839
rect 1741 784 1745 827
rect 1775 802 1779 876
rect 1767 790 1779 802
rect 1845 833 1849 916
rect 1905 839 1909 916
rect 1845 821 1854 833
rect 1906 827 1909 839
rect 1761 784 1765 790
rect 1845 764 1849 821
rect 1903 811 1909 827
rect 1925 839 1929 916
rect 1925 827 1934 839
rect 1971 833 1975 916
rect 2045 873 2049 916
rect 2065 904 2069 916
rect 2085 908 2089 916
rect 2085 904 2100 908
rect 2065 900 2080 904
rect 2074 893 2080 900
rect 2045 861 2053 873
rect 2065 861 2072 873
rect 1925 811 1931 827
rect 1966 821 1975 833
rect 1903 804 1917 811
rect 1913 784 1917 804
rect 1923 804 1931 811
rect 1923 784 1927 804
rect 1971 764 1975 821
rect 2068 804 2072 861
rect 2076 804 2080 881
rect 2094 873 2100 904
rect 2084 861 2094 873
rect 2084 804 2088 861
rect 2131 833 2135 916
rect 2196 872 2200 876
rect 2182 864 2200 872
rect 2182 853 2186 864
rect 2126 821 2135 833
rect 2131 764 2135 821
rect 2182 796 2186 841
rect 2204 819 2208 876
rect 2226 873 2230 916
rect 2226 861 2233 873
rect 2206 807 2215 819
rect 2182 789 2195 796
rect 2191 784 2195 789
rect 2211 784 2215 807
rect 2231 784 2235 861
rect 2305 819 2309 876
rect 2325 862 2329 876
rect 2345 862 2349 876
rect 2325 856 2340 862
rect 2345 856 2361 862
rect 2334 833 2340 856
rect 2305 807 2314 819
rect 2312 764 2316 807
rect 2334 784 2338 821
rect 2354 819 2361 856
rect 2391 833 2395 916
rect 2451 908 2455 916
rect 2440 904 2455 908
rect 2471 904 2475 916
rect 2440 873 2446 904
rect 2460 900 2475 904
rect 2460 893 2466 900
rect 2446 861 2456 873
rect 2386 821 2395 833
rect 2354 794 2361 807
rect 2342 788 2361 794
rect 2342 784 2346 788
rect 2391 764 2395 821
rect 2452 804 2456 861
rect 2460 804 2464 881
rect 2491 873 2495 916
rect 2468 861 2475 873
rect 2487 861 2495 873
rect 2565 873 2569 916
rect 2585 904 2589 916
rect 2605 908 2609 916
rect 2605 904 2620 908
rect 2585 900 2600 904
rect 2594 893 2600 900
rect 2565 861 2573 873
rect 2585 861 2592 873
rect 2468 804 2472 861
rect 2588 804 2592 861
rect 2596 804 2600 881
rect 2614 873 2620 904
rect 2604 861 2614 873
rect 2651 862 2655 876
rect 2671 862 2675 876
rect 2604 804 2608 861
rect 2639 856 2655 862
rect 2660 856 2675 862
rect 2639 819 2646 856
rect 2660 833 2666 856
rect 2639 794 2646 807
rect 2639 788 2658 794
rect 2654 784 2658 788
rect 2662 784 2666 821
rect 2691 819 2695 876
rect 2765 839 2769 916
rect 2766 827 2769 839
rect 2686 807 2695 819
rect 2763 811 2769 827
rect 2785 839 2789 916
rect 2855 872 2859 876
rect 2845 868 2859 872
rect 2845 853 2849 868
rect 2847 841 2849 853
rect 2785 827 2794 839
rect 2785 811 2791 827
rect 2684 764 2688 807
rect 2763 804 2777 811
rect 2773 784 2777 804
rect 2783 804 2791 811
rect 2783 784 2787 804
rect 2845 784 2849 841
rect 2865 819 2869 876
rect 2895 872 2899 876
rect 2885 868 2899 872
rect 2905 872 2909 876
rect 2905 868 2919 872
rect 2885 819 2891 868
rect 2914 853 2919 868
rect 2885 807 2894 819
rect 2865 784 2869 807
rect 2885 784 2889 807
rect 2914 795 2920 841
rect 2905 791 2920 795
rect 2965 833 2969 916
rect 3037 853 3041 876
rect 3026 841 3041 853
rect 3045 853 3049 876
rect 3117 853 3121 876
rect 3045 841 3054 853
rect 3106 841 3121 853
rect 3125 853 3129 876
rect 3125 841 3134 853
rect 2965 821 2974 833
rect 2905 784 2909 791
rect 2965 764 2969 821
rect 3025 764 3029 841
rect 3045 764 3049 841
rect 3105 764 3109 841
rect 3125 764 3129 841
rect 3171 833 3175 916
rect 3236 872 3240 876
rect 3222 864 3240 872
rect 3222 853 3226 864
rect 3166 821 3175 833
rect 3171 764 3175 821
rect 3222 796 3226 841
rect 3244 819 3248 876
rect 3266 873 3270 916
rect 3266 861 3273 873
rect 3246 807 3255 819
rect 3222 789 3235 796
rect 3231 784 3235 789
rect 3251 784 3255 807
rect 3271 784 3275 861
rect 3331 839 3335 916
rect 3326 827 3335 839
rect 3329 811 3335 827
rect 3351 839 3355 916
rect 3433 913 3437 936
rect 3429 906 3437 913
rect 3429 877 3433 906
rect 3441 896 3445 936
rect 3461 884 3465 916
rect 3469 912 3473 916
rect 3469 910 3505 912
rect 3469 908 3493 910
rect 3411 864 3415 876
rect 3429 871 3437 877
rect 3411 852 3413 864
rect 3351 827 3354 839
rect 3351 811 3357 827
rect 3329 804 3337 811
rect 3333 784 3337 804
rect 3343 804 3357 811
rect 3343 784 3347 804
rect 3411 784 3415 852
rect 3433 825 3437 871
rect 3433 764 3437 813
rect 3461 789 3467 884
rect 3443 785 3467 789
rect 3443 764 3447 785
rect 3463 780 3481 781
rect 3463 776 3493 780
rect 3463 764 3467 776
rect 3501 772 3505 898
rect 3515 890 3519 916
rect 3535 910 3539 916
rect 3471 768 3505 772
rect 3471 764 3475 768
rect 3517 764 3521 878
rect 3533 788 3537 898
rect 3547 876 3551 916
rect 3542 864 3545 876
rect 3542 800 3546 864
rect 3567 857 3571 916
rect 3562 849 3571 857
rect 3562 820 3566 849
rect 3581 834 3585 916
rect 3601 833 3605 876
rect 3651 853 3655 916
rect 3673 870 3677 876
rect 3675 858 3677 870
rect 3646 841 3655 853
rect 3542 796 3575 800
rect 3541 776 3543 788
rect 3539 764 3543 776
rect 3549 776 3551 788
rect 3549 764 3553 776
rect 3571 764 3575 796
rect 3581 764 3585 822
rect 3601 784 3605 821
rect 3651 764 3655 841
rect 3735 833 3739 876
rect 3755 834 3759 916
rect 3769 857 3773 916
rect 3789 876 3793 916
rect 3801 910 3805 916
rect 3795 864 3798 876
rect 3769 849 3778 857
rect 3675 790 3677 802
rect 3673 784 3677 790
rect 3735 784 3739 821
rect 3755 764 3759 822
rect 3774 820 3778 849
rect 3794 800 3798 864
rect 3765 796 3798 800
rect 3765 764 3769 796
rect 3803 788 3807 898
rect 3821 890 3825 916
rect 3867 912 3871 916
rect 3835 910 3871 912
rect 3847 908 3871 910
rect 3789 776 3791 788
rect 3787 764 3791 776
rect 3797 776 3799 788
rect 3797 764 3801 776
rect 3819 764 3823 878
rect 3835 772 3839 898
rect 3875 884 3879 916
rect 3895 896 3899 936
rect 3903 913 3907 936
rect 3903 906 3911 913
rect 3873 789 3879 884
rect 3907 877 3911 906
rect 3903 871 3911 877
rect 3903 825 3907 871
rect 3925 864 3929 876
rect 3990 873 3994 916
rect 4093 913 4097 936
rect 4089 906 4097 913
rect 4089 877 4093 906
rect 4101 896 4105 936
rect 4121 884 4125 916
rect 4129 912 4133 916
rect 4129 910 4165 912
rect 4129 908 4153 910
rect 3927 852 3929 864
rect 3987 861 3994 873
rect 3873 785 3897 789
rect 3859 780 3877 781
rect 3847 776 3877 780
rect 3835 768 3869 772
rect 3865 764 3869 768
rect 3873 764 3877 776
rect 3893 764 3897 785
rect 3903 764 3907 813
rect 3925 784 3929 852
rect 3985 784 3989 861
rect 4012 819 4016 876
rect 4020 872 4024 876
rect 4020 864 4038 872
rect 4034 853 4038 864
rect 4071 864 4075 876
rect 4089 871 4097 877
rect 4071 852 4073 864
rect 4005 807 4014 819
rect 4005 784 4009 807
rect 4034 796 4038 841
rect 4025 789 4038 796
rect 4025 784 4029 789
rect 4071 784 4075 852
rect 4093 825 4097 871
rect 4093 764 4097 813
rect 4121 789 4127 884
rect 4103 785 4127 789
rect 4103 764 4107 785
rect 4123 780 4141 781
rect 4123 776 4153 780
rect 4123 764 4127 776
rect 4161 772 4165 898
rect 4175 890 4179 916
rect 4195 910 4199 916
rect 4131 768 4165 772
rect 4131 764 4135 768
rect 4177 764 4181 878
rect 4193 788 4197 898
rect 4207 876 4211 916
rect 4202 864 4205 876
rect 4202 800 4206 864
rect 4227 857 4231 916
rect 4222 849 4231 857
rect 4222 820 4226 849
rect 4241 834 4245 916
rect 4261 833 4265 876
rect 4315 833 4319 876
rect 4335 834 4339 916
rect 4349 857 4353 916
rect 4369 876 4373 916
rect 4381 910 4385 916
rect 4375 864 4378 876
rect 4349 849 4358 857
rect 4202 796 4235 800
rect 4201 776 4203 788
rect 4199 764 4203 776
rect 4209 776 4211 788
rect 4209 764 4213 776
rect 4231 764 4235 796
rect 4241 764 4245 822
rect 4261 784 4265 821
rect 4315 784 4319 821
rect 4335 764 4339 822
rect 4354 820 4358 849
rect 4374 800 4378 864
rect 4345 796 4378 800
rect 4345 764 4349 796
rect 4383 788 4387 898
rect 4401 890 4405 916
rect 4447 912 4451 916
rect 4415 910 4451 912
rect 4427 908 4451 910
rect 4369 776 4371 788
rect 4367 764 4371 776
rect 4377 776 4379 788
rect 4377 764 4381 776
rect 4399 764 4403 878
rect 4415 772 4419 898
rect 4455 884 4459 916
rect 4475 896 4479 936
rect 4483 913 4487 936
rect 4483 906 4491 913
rect 4453 789 4459 884
rect 4487 877 4491 906
rect 4483 871 4491 877
rect 4483 825 4487 871
rect 4505 864 4509 876
rect 4556 872 4560 876
rect 4507 852 4509 864
rect 4542 864 4560 872
rect 4542 853 4546 864
rect 4453 785 4477 789
rect 4439 780 4457 781
rect 4427 776 4457 780
rect 4415 768 4449 772
rect 4445 764 4449 768
rect 4453 764 4457 776
rect 4473 764 4477 785
rect 4483 764 4487 813
rect 4505 784 4509 852
rect 4542 796 4546 841
rect 4564 819 4568 876
rect 4586 873 4590 916
rect 4586 861 4593 873
rect 4656 872 4660 876
rect 4642 864 4660 872
rect 4566 807 4575 819
rect 4542 789 4555 796
rect 4551 784 4555 789
rect 4571 784 4575 807
rect 4591 784 4595 861
rect 4642 853 4646 864
rect 4642 796 4646 841
rect 4664 819 4668 876
rect 4686 873 4690 916
rect 4686 861 4693 873
rect 4666 807 4675 819
rect 4642 789 4655 796
rect 4651 784 4655 789
rect 4671 784 4675 807
rect 4691 784 4695 861
rect 53 740 57 744
rect 63 740 67 744
rect 135 740 139 744
rect 155 740 159 744
rect 165 740 169 744
rect 225 740 229 744
rect 245 740 249 744
rect 265 740 269 744
rect 346 740 350 744
rect 354 740 358 744
rect 374 740 378 744
rect 382 740 386 744
rect 443 740 447 744
rect 465 740 469 744
rect 511 740 515 744
rect 585 740 589 744
rect 652 740 656 744
rect 674 740 678 744
rect 682 740 686 744
rect 732 740 736 744
rect 740 740 744 744
rect 748 740 752 744
rect 855 740 859 744
rect 875 740 879 744
rect 885 740 889 744
rect 933 740 937 744
rect 943 740 947 744
rect 1048 740 1052 744
rect 1056 740 1060 744
rect 1064 740 1068 744
rect 1111 740 1115 744
rect 1131 740 1135 744
rect 1151 740 1155 744
rect 1248 740 1252 744
rect 1256 740 1260 744
rect 1264 740 1268 744
rect 1311 740 1315 744
rect 1371 740 1375 744
rect 1391 740 1395 744
rect 1411 740 1415 744
rect 1493 740 1497 744
rect 1503 740 1507 744
rect 1553 740 1557 744
rect 1563 740 1567 744
rect 1645 740 1649 744
rect 1665 740 1669 744
rect 1685 740 1689 744
rect 1731 740 1735 744
rect 1741 740 1745 744
rect 1761 740 1765 744
rect 1845 740 1849 744
rect 1913 740 1917 744
rect 1923 740 1927 744
rect 1971 740 1975 744
rect 2068 740 2072 744
rect 2076 740 2080 744
rect 2084 740 2088 744
rect 2131 740 2135 744
rect 2191 740 2195 744
rect 2211 740 2215 744
rect 2231 740 2235 744
rect 2312 740 2316 744
rect 2334 740 2338 744
rect 2342 740 2346 744
rect 2391 740 2395 744
rect 2452 740 2456 744
rect 2460 740 2464 744
rect 2468 740 2472 744
rect 2588 740 2592 744
rect 2596 740 2600 744
rect 2604 740 2608 744
rect 2654 740 2658 744
rect 2662 740 2666 744
rect 2684 740 2688 744
rect 2773 740 2777 744
rect 2783 740 2787 744
rect 2845 740 2849 744
rect 2865 740 2869 744
rect 2885 740 2889 744
rect 2905 740 2909 744
rect 2965 740 2969 744
rect 3025 740 3029 744
rect 3045 740 3049 744
rect 3105 740 3109 744
rect 3125 740 3129 744
rect 3171 740 3175 744
rect 3231 740 3235 744
rect 3251 740 3255 744
rect 3271 740 3275 744
rect 3333 740 3337 744
rect 3343 740 3347 744
rect 3411 740 3415 744
rect 3433 740 3437 744
rect 3443 740 3447 744
rect 3463 740 3467 744
rect 3471 740 3475 744
rect 3517 740 3521 744
rect 3539 740 3543 744
rect 3549 740 3553 744
rect 3571 740 3575 744
rect 3581 740 3585 744
rect 3601 740 3605 744
rect 3651 740 3655 744
rect 3673 740 3677 744
rect 3735 740 3739 744
rect 3755 740 3759 744
rect 3765 740 3769 744
rect 3787 740 3791 744
rect 3797 740 3801 744
rect 3819 740 3823 744
rect 3865 740 3869 744
rect 3873 740 3877 744
rect 3893 740 3897 744
rect 3903 740 3907 744
rect 3925 740 3929 744
rect 3985 740 3989 744
rect 4005 740 4009 744
rect 4025 740 4029 744
rect 4071 740 4075 744
rect 4093 740 4097 744
rect 4103 740 4107 744
rect 4123 740 4127 744
rect 4131 740 4135 744
rect 4177 740 4181 744
rect 4199 740 4203 744
rect 4209 740 4213 744
rect 4231 740 4235 744
rect 4241 740 4245 744
rect 4261 740 4265 744
rect 4315 740 4319 744
rect 4335 740 4339 744
rect 4345 740 4349 744
rect 4367 740 4371 744
rect 4377 740 4381 744
rect 4399 740 4403 744
rect 4445 740 4449 744
rect 4453 740 4457 744
rect 4473 740 4477 744
rect 4483 740 4487 744
rect 4505 740 4509 744
rect 4551 740 4555 744
rect 4571 740 4575 744
rect 4591 740 4595 744
rect 4651 740 4655 744
rect 4671 740 4675 744
rect 4691 740 4695 744
rect 45 716 49 720
rect 65 716 69 720
rect 132 716 136 720
rect 154 716 158 720
rect 162 716 166 720
rect 211 716 215 720
rect 292 716 296 720
rect 314 716 318 720
rect 322 716 326 720
rect 372 716 376 720
rect 380 716 384 720
rect 388 716 392 720
rect 485 716 489 720
rect 505 716 509 720
rect 525 716 529 720
rect 583 716 587 720
rect 605 716 609 720
rect 665 716 669 720
rect 685 716 689 720
rect 705 716 709 720
rect 763 716 767 720
rect 785 716 789 720
rect 831 716 835 720
rect 841 716 845 720
rect 861 716 865 720
rect 931 716 935 720
rect 951 716 955 720
rect 971 716 975 720
rect 1045 716 1049 720
rect 1065 716 1069 720
rect 1085 716 1089 720
rect 1145 716 1149 720
rect 1194 716 1198 720
rect 1202 716 1206 720
rect 1224 716 1228 720
rect 1305 716 1309 720
rect 1351 716 1355 720
rect 1371 716 1375 720
rect 1391 716 1395 720
rect 1451 716 1455 720
rect 1471 716 1475 720
rect 1491 716 1495 720
rect 1572 716 1576 720
rect 1594 716 1598 720
rect 1602 716 1606 720
rect 1654 716 1658 720
rect 1662 716 1666 720
rect 1684 716 1688 720
rect 1752 716 1756 720
rect 1760 716 1764 720
rect 1768 716 1772 720
rect 1851 716 1855 720
rect 1871 716 1875 720
rect 1891 716 1895 720
rect 1972 716 1976 720
rect 1994 716 1998 720
rect 2002 716 2006 720
rect 2051 716 2055 720
rect 2071 716 2075 720
rect 2091 716 2095 720
rect 2188 716 2192 720
rect 2196 716 2200 720
rect 2204 716 2208 720
rect 2265 716 2269 720
rect 2285 716 2289 720
rect 2305 716 2309 720
rect 2351 716 2355 720
rect 2371 716 2375 720
rect 2391 716 2395 720
rect 2452 716 2456 720
rect 2460 716 2464 720
rect 2468 716 2472 720
rect 2552 716 2556 720
rect 2560 716 2564 720
rect 2568 716 2572 720
rect 2665 716 2669 720
rect 2712 716 2716 720
rect 2720 716 2724 720
rect 2728 716 2732 720
rect 2815 716 2819 720
rect 2835 716 2839 720
rect 2845 716 2849 720
rect 2867 716 2871 720
rect 2877 716 2881 720
rect 2899 716 2903 720
rect 2945 716 2949 720
rect 2953 716 2957 720
rect 2973 716 2977 720
rect 2983 716 2987 720
rect 3005 716 3009 720
rect 3051 716 3055 720
rect 3071 716 3075 720
rect 3091 716 3095 720
rect 3151 716 3155 720
rect 3211 716 3215 720
rect 3272 716 3276 720
rect 3280 716 3284 720
rect 3288 716 3292 720
rect 3385 716 3389 720
rect 3453 716 3457 720
rect 3463 716 3467 720
rect 3525 716 3529 720
rect 3545 716 3549 720
rect 3565 716 3569 720
rect 3615 716 3619 720
rect 3635 716 3639 720
rect 3645 716 3649 720
rect 3667 716 3671 720
rect 3677 716 3681 720
rect 3699 716 3703 720
rect 3745 716 3749 720
rect 3753 716 3757 720
rect 3773 716 3777 720
rect 3783 716 3787 720
rect 3805 716 3809 720
rect 3851 716 3855 720
rect 3871 716 3875 720
rect 3891 716 3895 720
rect 3973 716 3977 720
rect 3983 716 3987 720
rect 4031 716 4035 720
rect 4053 716 4057 720
rect 4063 716 4067 720
rect 4083 716 4087 720
rect 4091 716 4095 720
rect 4137 716 4141 720
rect 4159 716 4163 720
rect 4169 716 4173 720
rect 4191 716 4195 720
rect 4201 716 4205 720
rect 4221 716 4225 720
rect 4273 716 4277 720
rect 4283 716 4287 720
rect 4353 716 4357 720
rect 4363 716 4367 720
rect 4445 716 4449 720
rect 4465 716 4469 720
rect 4485 716 4489 720
rect 4535 716 4539 720
rect 4555 716 4559 720
rect 4565 716 4569 720
rect 4587 716 4591 720
rect 4597 716 4601 720
rect 4619 716 4623 720
rect 4665 716 4669 720
rect 4673 716 4677 720
rect 4693 716 4697 720
rect 4703 716 4707 720
rect 4725 716 4729 720
rect 45 619 49 696
rect 65 619 69 696
rect 132 653 136 696
rect 125 641 134 653
rect 46 607 61 619
rect 57 584 61 607
rect 65 607 74 619
rect 65 584 69 607
rect 125 584 129 641
rect 154 639 158 676
rect 162 672 166 676
rect 162 666 181 672
rect 174 653 181 666
rect 154 604 160 627
rect 174 604 181 641
rect 211 639 215 696
rect 292 653 296 696
rect 206 627 215 639
rect 145 598 160 604
rect 165 598 181 604
rect 145 584 149 598
rect 165 584 169 598
rect 211 544 215 627
rect 285 641 294 653
rect 285 584 289 641
rect 314 639 318 676
rect 322 672 326 676
rect 322 666 341 672
rect 334 653 341 666
rect 314 604 320 627
rect 334 604 341 641
rect 305 598 320 604
rect 325 598 341 604
rect 372 599 376 656
rect 305 584 309 598
rect 325 584 329 598
rect 366 587 376 599
rect 360 556 366 587
rect 380 579 384 656
rect 388 599 392 656
rect 485 599 489 676
rect 505 653 509 676
rect 525 671 529 676
rect 525 664 538 671
rect 505 641 514 653
rect 388 587 395 599
rect 407 587 415 599
rect 487 587 494 599
rect 380 560 386 567
rect 380 556 395 560
rect 360 552 375 556
rect 371 544 375 552
rect 391 544 395 556
rect 411 544 415 587
rect 490 544 494 587
rect 512 584 516 641
rect 534 619 538 664
rect 583 670 587 676
rect 583 658 585 670
rect 605 619 609 696
rect 605 607 614 619
rect 534 596 538 607
rect 520 588 538 596
rect 583 590 585 602
rect 520 584 524 588
rect 583 584 587 590
rect 605 544 609 607
rect 665 599 669 676
rect 685 653 689 676
rect 705 671 709 676
rect 705 664 718 671
rect 685 641 694 653
rect 667 587 674 599
rect 670 544 674 587
rect 692 584 696 641
rect 714 619 718 664
rect 763 670 767 676
rect 763 658 765 670
rect 785 619 789 696
rect 831 619 835 676
rect 841 633 845 676
rect 861 670 865 676
rect 931 671 935 676
rect 867 658 879 670
rect 841 621 854 633
rect 785 607 794 619
rect 826 607 835 619
rect 714 596 718 607
rect 700 588 718 596
rect 763 590 765 602
rect 700 584 704 588
rect 763 584 767 590
rect 785 544 789 607
rect 831 544 835 607
rect 853 544 857 621
rect 875 584 879 658
rect 922 664 935 671
rect 922 619 926 664
rect 951 653 955 676
rect 946 641 955 653
rect 922 596 926 607
rect 922 588 940 596
rect 936 584 940 588
rect 944 584 948 641
rect 971 599 975 676
rect 1045 599 1049 676
rect 1065 653 1069 676
rect 1085 671 1089 676
rect 1085 664 1098 671
rect 1065 641 1074 653
rect 966 587 973 599
rect 1047 587 1054 599
rect 966 544 970 587
rect 1050 544 1054 587
rect 1072 584 1076 641
rect 1094 619 1098 664
rect 1145 653 1149 676
rect 1194 672 1198 676
rect 1179 666 1198 672
rect 1179 653 1186 666
rect 1145 641 1154 653
rect 1094 596 1098 607
rect 1080 588 1098 596
rect 1080 584 1084 588
rect 1145 584 1149 641
rect 1179 604 1186 641
rect 1202 639 1206 676
rect 1224 653 1228 696
rect 1226 641 1235 653
rect 1200 604 1206 627
rect 1179 598 1195 604
rect 1200 598 1215 604
rect 1191 584 1195 598
rect 1211 584 1215 598
rect 1231 584 1235 641
rect 1305 639 1309 696
rect 1351 671 1355 676
rect 1342 664 1355 671
rect 1305 627 1314 639
rect 1305 544 1309 627
rect 1342 619 1346 664
rect 1371 653 1375 676
rect 1366 641 1375 653
rect 1342 596 1346 607
rect 1342 588 1360 596
rect 1356 584 1360 588
rect 1364 584 1368 641
rect 1391 599 1395 676
rect 1451 671 1455 676
rect 1442 664 1455 671
rect 1442 619 1446 664
rect 1471 653 1475 676
rect 1466 641 1475 653
rect 1386 587 1393 599
rect 1442 596 1446 607
rect 1442 588 1460 596
rect 1386 544 1390 587
rect 1456 584 1460 588
rect 1464 584 1468 641
rect 1491 599 1495 676
rect 1572 653 1576 696
rect 1565 641 1574 653
rect 1486 587 1493 599
rect 1486 544 1490 587
rect 1565 584 1569 641
rect 1594 639 1598 676
rect 1602 672 1606 676
rect 1654 672 1658 676
rect 1602 666 1621 672
rect 1614 653 1621 666
rect 1639 666 1658 672
rect 1639 653 1646 666
rect 1594 604 1600 627
rect 1614 604 1621 641
rect 1585 598 1600 604
rect 1605 598 1621 604
rect 1639 604 1646 641
rect 1662 639 1666 676
rect 1684 653 1688 696
rect 1851 671 1855 676
rect 1842 664 1855 671
rect 1686 641 1695 653
rect 1660 604 1666 627
rect 1639 598 1655 604
rect 1660 598 1675 604
rect 1585 584 1589 598
rect 1605 584 1609 598
rect 1651 584 1655 598
rect 1671 584 1675 598
rect 1691 584 1695 641
rect 1752 599 1756 656
rect 1746 587 1756 599
rect 1740 556 1746 587
rect 1760 579 1764 656
rect 1768 599 1772 656
rect 1842 619 1846 664
rect 1871 653 1875 676
rect 1866 641 1875 653
rect 1768 587 1775 599
rect 1787 587 1795 599
rect 1842 596 1846 607
rect 1842 588 1860 596
rect 1760 560 1766 567
rect 1760 556 1775 560
rect 1740 552 1755 556
rect 1751 544 1755 552
rect 1771 544 1775 556
rect 1791 544 1795 587
rect 1856 584 1860 588
rect 1864 584 1868 641
rect 1891 599 1895 676
rect 1972 653 1976 696
rect 1965 641 1974 653
rect 1886 587 1893 599
rect 1886 544 1890 587
rect 1965 584 1969 641
rect 1994 639 1998 676
rect 2002 672 2006 676
rect 2002 666 2021 672
rect 2051 671 2055 676
rect 2014 653 2021 666
rect 2042 664 2055 671
rect 1994 604 2000 627
rect 2014 604 2021 641
rect 2042 619 2046 664
rect 2071 653 2075 676
rect 2066 641 2075 653
rect 1985 598 2000 604
rect 2005 598 2021 604
rect 1985 584 1989 598
rect 2005 584 2009 598
rect 2042 596 2046 607
rect 2042 588 2060 596
rect 2056 584 2060 588
rect 2064 584 2068 641
rect 2091 599 2095 676
rect 2188 599 2192 656
rect 2086 587 2093 599
rect 2165 587 2173 599
rect 2185 587 2192 599
rect 2086 544 2090 587
rect 2165 544 2169 587
rect 2196 579 2200 656
rect 2204 599 2208 656
rect 2265 599 2269 676
rect 2285 653 2289 676
rect 2305 671 2309 676
rect 2351 671 2355 676
rect 2305 664 2318 671
rect 2285 641 2294 653
rect 2204 587 2214 599
rect 2267 587 2274 599
rect 2194 560 2200 567
rect 2185 556 2200 560
rect 2214 556 2220 587
rect 2185 544 2189 556
rect 2205 552 2220 556
rect 2205 544 2209 552
rect 2270 544 2274 587
rect 2292 584 2296 641
rect 2314 619 2318 664
rect 2342 664 2355 671
rect 2342 619 2346 664
rect 2371 653 2375 676
rect 2366 641 2375 653
rect 2314 596 2318 607
rect 2300 588 2318 596
rect 2342 596 2346 607
rect 2342 588 2360 596
rect 2300 584 2304 588
rect 2356 584 2360 588
rect 2364 584 2368 641
rect 2391 599 2395 676
rect 2452 599 2456 656
rect 2386 587 2393 599
rect 2446 587 2456 599
rect 2386 544 2390 587
rect 2440 556 2446 587
rect 2460 579 2464 656
rect 2468 599 2472 656
rect 2552 599 2556 656
rect 2468 587 2475 599
rect 2487 587 2495 599
rect 2546 587 2556 599
rect 2460 560 2466 567
rect 2460 556 2475 560
rect 2440 552 2455 556
rect 2451 544 2455 552
rect 2471 544 2475 556
rect 2491 544 2495 587
rect 2540 556 2546 587
rect 2560 579 2564 656
rect 2568 599 2572 656
rect 2665 639 2669 696
rect 2665 627 2674 639
rect 2568 587 2575 599
rect 2587 587 2595 599
rect 2560 560 2566 567
rect 2560 556 2575 560
rect 2540 552 2555 556
rect 2551 544 2555 552
rect 2571 544 2575 556
rect 2591 544 2595 587
rect 2665 544 2669 627
rect 2712 599 2716 656
rect 2706 587 2716 599
rect 2700 556 2706 587
rect 2720 579 2724 656
rect 2728 599 2732 656
rect 2815 639 2819 676
rect 2835 638 2839 696
rect 2845 664 2849 696
rect 2867 684 2871 696
rect 2869 672 2871 684
rect 2877 684 2881 696
rect 2877 672 2879 684
rect 2845 660 2878 664
rect 2728 587 2735 599
rect 2747 587 2755 599
rect 2720 560 2726 567
rect 2720 556 2735 560
rect 2700 552 2715 556
rect 2711 544 2715 552
rect 2731 544 2735 556
rect 2751 544 2755 587
rect 2815 584 2819 627
rect 2835 544 2839 626
rect 2854 611 2858 640
rect 2849 603 2858 611
rect 2849 544 2853 603
rect 2874 596 2878 660
rect 2875 584 2878 596
rect 2869 544 2873 584
rect 2883 562 2887 672
rect 2899 582 2903 696
rect 2945 692 2949 696
rect 2915 688 2949 692
rect 2881 544 2885 550
rect 2901 544 2905 570
rect 2915 562 2919 688
rect 2953 684 2957 696
rect 2927 680 2957 684
rect 2939 679 2957 680
rect 2973 675 2977 696
rect 2953 671 2977 675
rect 2953 576 2959 671
rect 2983 647 2987 696
rect 2983 589 2987 635
rect 3005 608 3009 676
rect 3051 671 3055 676
rect 3042 664 3055 671
rect 3042 619 3046 664
rect 3071 653 3075 676
rect 3066 641 3075 653
rect 3007 596 3009 608
rect 2983 583 2991 589
rect 3005 584 3009 596
rect 3042 596 3046 607
rect 3042 588 3060 596
rect 3056 584 3060 588
rect 3064 584 3068 641
rect 3091 599 3095 676
rect 3151 639 3155 696
rect 3211 639 3215 696
rect 3146 627 3155 639
rect 3206 627 3215 639
rect 3086 587 3093 599
rect 2927 550 2951 552
rect 2915 548 2951 550
rect 2947 544 2951 548
rect 2955 544 2959 576
rect 2975 524 2979 564
rect 2987 554 2991 583
rect 2983 547 2991 554
rect 2983 524 2987 547
rect 3086 544 3090 587
rect 3151 544 3155 627
rect 3211 544 3215 627
rect 3272 599 3276 656
rect 3266 587 3276 599
rect 3260 556 3266 587
rect 3280 579 3284 656
rect 3288 599 3292 656
rect 3385 639 3389 696
rect 3453 656 3457 676
rect 3443 649 3457 656
rect 3463 656 3467 676
rect 3463 649 3471 656
rect 3385 627 3394 639
rect 3443 633 3449 649
rect 3288 587 3295 599
rect 3307 587 3315 599
rect 3280 560 3286 567
rect 3280 556 3295 560
rect 3260 552 3275 556
rect 3271 544 3275 552
rect 3291 544 3295 556
rect 3311 544 3315 587
rect 3385 544 3389 627
rect 3446 621 3449 633
rect 3445 544 3449 621
rect 3465 633 3471 649
rect 3465 621 3474 633
rect 3465 544 3469 621
rect 3525 599 3529 676
rect 3545 653 3549 676
rect 3565 671 3569 676
rect 3565 664 3578 671
rect 3545 641 3554 653
rect 3527 587 3534 599
rect 3530 544 3534 587
rect 3552 584 3556 641
rect 3574 619 3578 664
rect 3615 639 3619 676
rect 3635 638 3639 696
rect 3645 664 3649 696
rect 3667 684 3671 696
rect 3669 672 3671 684
rect 3677 684 3681 696
rect 3677 672 3679 684
rect 3645 660 3678 664
rect 3574 596 3578 607
rect 3560 588 3578 596
rect 3560 584 3564 588
rect 3615 584 3619 627
rect 3635 544 3639 626
rect 3654 611 3658 640
rect 3649 603 3658 611
rect 3649 544 3653 603
rect 3674 596 3678 660
rect 3675 584 3678 596
rect 3669 544 3673 584
rect 3683 562 3687 672
rect 3699 582 3703 696
rect 3745 692 3749 696
rect 3715 688 3749 692
rect 3681 544 3685 550
rect 3701 544 3705 570
rect 3715 562 3719 688
rect 3753 684 3757 696
rect 3727 680 3757 684
rect 3739 679 3757 680
rect 3773 675 3777 696
rect 3753 671 3777 675
rect 3753 576 3759 671
rect 3783 647 3787 696
rect 3783 589 3787 635
rect 3805 608 3809 676
rect 3851 671 3855 676
rect 3842 664 3855 671
rect 3842 619 3846 664
rect 3871 653 3875 676
rect 3866 641 3875 653
rect 3807 596 3809 608
rect 3783 583 3791 589
rect 3805 584 3809 596
rect 3842 596 3846 607
rect 3842 588 3860 596
rect 3856 584 3860 588
rect 3864 584 3868 641
rect 3891 599 3895 676
rect 3973 656 3977 676
rect 3963 649 3977 656
rect 3983 656 3987 676
rect 3983 649 3991 656
rect 3963 633 3969 649
rect 3966 621 3969 633
rect 3886 587 3893 599
rect 3727 550 3751 552
rect 3715 548 3751 550
rect 3747 544 3751 548
rect 3755 544 3759 576
rect 3775 524 3779 564
rect 3787 554 3791 583
rect 3783 547 3791 554
rect 3783 524 3787 547
rect 3886 544 3890 587
rect 3965 544 3969 621
rect 3985 633 3991 649
rect 3985 621 3994 633
rect 3985 544 3989 621
rect 4031 608 4035 676
rect 4053 647 4057 696
rect 4063 675 4067 696
rect 4083 684 4087 696
rect 4091 692 4095 696
rect 4091 688 4125 692
rect 4083 680 4113 684
rect 4083 679 4101 680
rect 4063 671 4087 675
rect 4031 596 4033 608
rect 4031 584 4035 596
rect 4053 589 4057 635
rect 4049 583 4057 589
rect 4049 554 4053 583
rect 4081 576 4087 671
rect 4049 547 4057 554
rect 4053 524 4057 547
rect 4061 524 4065 564
rect 4081 544 4085 576
rect 4121 562 4125 688
rect 4137 582 4141 696
rect 4159 684 4163 696
rect 4161 672 4163 684
rect 4169 684 4173 696
rect 4169 672 4171 684
rect 4089 550 4113 552
rect 4089 548 4125 550
rect 4089 544 4093 548
rect 4135 544 4139 570
rect 4153 562 4157 672
rect 4191 664 4195 696
rect 4162 660 4195 664
rect 4162 596 4166 660
rect 4182 611 4186 640
rect 4201 638 4205 696
rect 4221 639 4225 676
rect 4273 656 4277 676
rect 4269 649 4277 656
rect 4283 656 4287 676
rect 4353 656 4357 676
rect 4283 649 4297 656
rect 4269 633 4275 649
rect 4182 603 4191 611
rect 4162 584 4165 596
rect 4155 544 4159 550
rect 4167 544 4171 584
rect 4187 544 4191 603
rect 4201 544 4205 626
rect 4221 584 4225 627
rect 4266 621 4275 633
rect 4271 544 4275 621
rect 4291 633 4297 649
rect 4349 649 4357 656
rect 4363 656 4367 676
rect 4363 649 4377 656
rect 4349 633 4355 649
rect 4291 621 4294 633
rect 4346 621 4355 633
rect 4291 544 4295 621
rect 4351 544 4355 621
rect 4371 633 4377 649
rect 4371 621 4374 633
rect 4371 544 4375 621
rect 4445 599 4449 676
rect 4465 653 4469 676
rect 4485 671 4489 676
rect 4485 664 4498 671
rect 4465 641 4474 653
rect 4447 587 4454 599
rect 4450 544 4454 587
rect 4472 584 4476 641
rect 4494 619 4498 664
rect 4535 639 4539 676
rect 4555 638 4559 696
rect 4565 664 4569 696
rect 4587 684 4591 696
rect 4589 672 4591 684
rect 4597 684 4601 696
rect 4597 672 4599 684
rect 4565 660 4598 664
rect 4494 596 4498 607
rect 4480 588 4498 596
rect 4480 584 4484 588
rect 4535 584 4539 627
rect 4555 544 4559 626
rect 4574 611 4578 640
rect 4569 603 4578 611
rect 4569 544 4573 603
rect 4594 596 4598 660
rect 4595 584 4598 596
rect 4589 544 4593 584
rect 4603 562 4607 672
rect 4619 582 4623 696
rect 4665 692 4669 696
rect 4635 688 4669 692
rect 4601 544 4605 550
rect 4621 544 4625 570
rect 4635 562 4639 688
rect 4673 684 4677 696
rect 4647 680 4677 684
rect 4659 679 4677 680
rect 4693 675 4697 696
rect 4673 671 4697 675
rect 4673 576 4679 671
rect 4703 647 4707 696
rect 4703 589 4707 635
rect 4725 608 4729 676
rect 4727 596 4729 608
rect 4703 583 4711 589
rect 4725 584 4729 596
rect 4647 550 4671 552
rect 4635 548 4671 550
rect 4667 544 4671 548
rect 4675 544 4679 576
rect 4695 524 4699 564
rect 4707 554 4711 583
rect 4703 547 4711 554
rect 4703 524 4707 547
rect 57 500 61 504
rect 65 500 69 504
rect 125 500 129 504
rect 145 500 149 504
rect 165 500 169 504
rect 211 500 215 504
rect 285 500 289 504
rect 305 500 309 504
rect 325 500 329 504
rect 371 500 375 504
rect 391 500 395 504
rect 411 500 415 504
rect 490 500 494 504
rect 512 500 516 504
rect 520 500 524 504
rect 583 500 587 504
rect 605 500 609 504
rect 670 500 674 504
rect 692 500 696 504
rect 700 500 704 504
rect 763 500 767 504
rect 785 500 789 504
rect 831 500 835 504
rect 853 500 857 504
rect 875 500 879 504
rect 936 500 940 504
rect 944 500 948 504
rect 966 500 970 504
rect 1050 500 1054 504
rect 1072 500 1076 504
rect 1080 500 1084 504
rect 1145 500 1149 504
rect 1191 500 1195 504
rect 1211 500 1215 504
rect 1231 500 1235 504
rect 1305 500 1309 504
rect 1356 500 1360 504
rect 1364 500 1368 504
rect 1386 500 1390 504
rect 1456 500 1460 504
rect 1464 500 1468 504
rect 1486 500 1490 504
rect 1565 500 1569 504
rect 1585 500 1589 504
rect 1605 500 1609 504
rect 1651 500 1655 504
rect 1671 500 1675 504
rect 1691 500 1695 504
rect 1751 500 1755 504
rect 1771 500 1775 504
rect 1791 500 1795 504
rect 1856 500 1860 504
rect 1864 500 1868 504
rect 1886 500 1890 504
rect 1965 500 1969 504
rect 1985 500 1989 504
rect 2005 500 2009 504
rect 2056 500 2060 504
rect 2064 500 2068 504
rect 2086 500 2090 504
rect 2165 500 2169 504
rect 2185 500 2189 504
rect 2205 500 2209 504
rect 2270 500 2274 504
rect 2292 500 2296 504
rect 2300 500 2304 504
rect 2356 500 2360 504
rect 2364 500 2368 504
rect 2386 500 2390 504
rect 2451 500 2455 504
rect 2471 500 2475 504
rect 2491 500 2495 504
rect 2551 500 2555 504
rect 2571 500 2575 504
rect 2591 500 2595 504
rect 2665 500 2669 504
rect 2711 500 2715 504
rect 2731 500 2735 504
rect 2751 500 2755 504
rect 2815 500 2819 504
rect 2835 500 2839 504
rect 2849 500 2853 504
rect 2869 500 2873 504
rect 2881 500 2885 504
rect 2901 500 2905 504
rect 2947 500 2951 504
rect 2955 500 2959 504
rect 2975 500 2979 504
rect 2983 500 2987 504
rect 3005 500 3009 504
rect 3056 500 3060 504
rect 3064 500 3068 504
rect 3086 500 3090 504
rect 3151 500 3155 504
rect 3211 500 3215 504
rect 3271 500 3275 504
rect 3291 500 3295 504
rect 3311 500 3315 504
rect 3385 500 3389 504
rect 3445 500 3449 504
rect 3465 500 3469 504
rect 3530 500 3534 504
rect 3552 500 3556 504
rect 3560 500 3564 504
rect 3615 500 3619 504
rect 3635 500 3639 504
rect 3649 500 3653 504
rect 3669 500 3673 504
rect 3681 500 3685 504
rect 3701 500 3705 504
rect 3747 500 3751 504
rect 3755 500 3759 504
rect 3775 500 3779 504
rect 3783 500 3787 504
rect 3805 500 3809 504
rect 3856 500 3860 504
rect 3864 500 3868 504
rect 3886 500 3890 504
rect 3965 500 3969 504
rect 3985 500 3989 504
rect 4031 500 4035 504
rect 4053 500 4057 504
rect 4061 500 4065 504
rect 4081 500 4085 504
rect 4089 500 4093 504
rect 4135 500 4139 504
rect 4155 500 4159 504
rect 4167 500 4171 504
rect 4187 500 4191 504
rect 4201 500 4205 504
rect 4221 500 4225 504
rect 4271 500 4275 504
rect 4291 500 4295 504
rect 4351 500 4355 504
rect 4371 500 4375 504
rect 4450 500 4454 504
rect 4472 500 4476 504
rect 4480 500 4484 504
rect 4535 500 4539 504
rect 4555 500 4559 504
rect 4569 500 4573 504
rect 4589 500 4593 504
rect 4601 500 4605 504
rect 4621 500 4625 504
rect 4667 500 4671 504
rect 4675 500 4679 504
rect 4695 500 4699 504
rect 4703 500 4707 504
rect 4725 500 4729 504
rect 31 476 35 480
rect 51 476 55 480
rect 111 476 115 480
rect 131 476 135 480
rect 205 476 209 480
rect 225 476 229 480
rect 285 476 289 480
rect 305 476 309 480
rect 361 476 365 480
rect 383 476 387 480
rect 405 476 409 480
rect 465 476 469 480
rect 485 476 489 480
rect 545 476 549 480
rect 565 476 569 480
rect 585 476 589 480
rect 645 476 649 480
rect 665 476 669 480
rect 685 476 689 480
rect 705 476 709 480
rect 777 476 781 480
rect 785 476 789 480
rect 845 476 849 480
rect 865 476 869 480
rect 911 476 915 480
rect 931 476 935 480
rect 1005 476 1009 480
rect 1025 476 1029 480
rect 1085 476 1089 480
rect 1105 476 1109 480
rect 1165 476 1169 480
rect 1185 476 1189 480
rect 1205 476 1209 480
rect 1225 476 1229 480
rect 1276 476 1280 480
rect 1284 476 1288 480
rect 1306 476 1310 480
rect 1397 476 1401 480
rect 1405 476 1409 480
rect 1456 476 1460 480
rect 1464 476 1468 480
rect 1486 476 1490 480
rect 1551 476 1555 480
rect 1625 476 1629 480
rect 1645 476 1649 480
rect 1665 476 1669 480
rect 1711 476 1715 480
rect 1771 476 1775 480
rect 1791 476 1795 480
rect 1811 476 1815 480
rect 1871 476 1875 480
rect 1891 476 1895 480
rect 1911 476 1915 480
rect 1971 476 1975 480
rect 1991 476 1995 480
rect 2051 476 2055 480
rect 2071 476 2075 480
rect 2131 476 2135 480
rect 2151 476 2155 480
rect 2237 476 2241 480
rect 2245 476 2249 480
rect 2305 476 2309 480
rect 2325 476 2329 480
rect 2371 476 2375 480
rect 2379 476 2383 480
rect 2451 476 2455 480
rect 2471 476 2475 480
rect 2491 476 2495 480
rect 2565 476 2569 480
rect 2625 476 2629 480
rect 2645 476 2649 480
rect 2665 476 2669 480
rect 2711 476 2715 480
rect 2731 476 2735 480
rect 2751 476 2755 480
rect 2811 476 2815 480
rect 2819 476 2823 480
rect 2905 476 2909 480
rect 2925 476 2929 480
rect 2990 476 2994 480
rect 3012 476 3016 480
rect 3020 476 3024 480
rect 3090 476 3094 480
rect 3112 476 3116 480
rect 3120 476 3124 480
rect 3197 476 3201 480
rect 3205 476 3209 480
rect 3265 476 3269 480
rect 3330 476 3334 480
rect 3352 476 3356 480
rect 3360 476 3364 480
rect 3425 476 3429 480
rect 3445 476 3449 480
rect 3465 476 3469 480
rect 3537 476 3541 480
rect 3545 476 3549 480
rect 3591 476 3595 480
rect 3601 476 3605 480
rect 3621 476 3625 480
rect 3691 476 3695 480
rect 3711 476 3715 480
rect 3771 476 3775 480
rect 3791 476 3795 480
rect 3870 476 3874 480
rect 3892 476 3896 480
rect 3900 476 3904 480
rect 3965 476 3969 480
rect 4025 476 4029 480
rect 4071 476 4075 480
rect 4093 476 4097 480
rect 4101 476 4105 480
rect 4121 476 4125 480
rect 4129 476 4133 480
rect 4175 476 4179 480
rect 4195 476 4199 480
rect 4207 476 4211 480
rect 4227 476 4231 480
rect 4241 476 4245 480
rect 4261 476 4265 480
rect 4325 476 4329 480
rect 4345 476 4349 480
rect 4410 476 4414 480
rect 4432 476 4436 480
rect 4440 476 4444 480
rect 4505 476 4509 480
rect 4551 476 4555 480
rect 4573 476 4577 480
rect 4581 476 4585 480
rect 4601 476 4605 480
rect 4609 476 4613 480
rect 4655 476 4659 480
rect 4675 476 4679 480
rect 4687 476 4691 480
rect 4707 476 4711 480
rect 4721 476 4725 480
rect 4741 476 4745 480
rect 31 359 35 436
rect 26 347 35 359
rect 29 331 35 347
rect 51 359 55 436
rect 111 359 115 436
rect 51 347 54 359
rect 106 347 115 359
rect 51 331 57 347
rect 29 324 37 331
rect 33 304 37 324
rect 43 324 57 331
rect 109 331 115 347
rect 131 359 135 436
rect 205 359 209 436
rect 131 347 134 359
rect 206 347 209 359
rect 131 331 137 347
rect 109 324 117 331
rect 43 304 47 324
rect 113 304 117 324
rect 123 324 137 331
rect 203 331 209 347
rect 225 359 229 436
rect 285 359 289 436
rect 225 347 234 359
rect 286 347 289 359
rect 225 331 231 347
rect 203 324 217 331
rect 123 304 127 324
rect 213 304 217 324
rect 223 324 231 331
rect 283 331 289 347
rect 305 359 309 436
rect 305 347 314 359
rect 305 331 311 347
rect 283 324 297 331
rect 223 304 227 324
rect 293 304 297 324
rect 303 324 311 331
rect 303 304 307 324
rect 361 322 365 396
rect 383 359 387 436
rect 405 373 409 436
rect 405 361 414 373
rect 386 347 399 359
rect 361 310 373 322
rect 375 304 379 310
rect 395 304 399 347
rect 405 304 409 361
rect 465 359 469 436
rect 466 347 469 359
rect 463 331 469 347
rect 485 359 489 436
rect 545 393 549 436
rect 565 424 569 436
rect 585 428 589 436
rect 585 424 600 428
rect 565 420 580 424
rect 574 413 580 420
rect 545 381 553 393
rect 565 381 572 393
rect 485 347 494 359
rect 485 331 491 347
rect 463 324 477 331
rect 473 304 477 324
rect 483 324 491 331
rect 568 324 572 381
rect 576 324 580 401
rect 594 393 600 424
rect 584 381 594 393
rect 584 324 588 381
rect 645 373 649 396
rect 646 361 649 373
rect 483 304 487 324
rect 640 313 646 361
rect 665 339 669 396
rect 685 374 689 396
rect 705 374 709 396
rect 685 368 698 374
rect 705 373 725 374
rect 777 373 781 396
rect 705 368 713 373
rect 694 339 698 368
rect 766 361 781 373
rect 785 373 789 396
rect 785 361 794 373
rect 667 327 669 339
rect 665 325 669 327
rect 665 318 678 325
rect 640 309 670 313
rect 666 304 670 309
rect 674 304 678 318
rect 694 304 698 327
rect 713 319 719 361
rect 702 312 719 319
rect 702 304 706 312
rect 765 284 769 361
rect 785 284 789 361
rect 845 359 849 436
rect 846 347 849 359
rect 843 331 849 347
rect 865 359 869 436
rect 911 359 915 436
rect 865 347 874 359
rect 906 347 915 359
rect 865 331 871 347
rect 843 324 857 331
rect 853 304 857 324
rect 863 324 871 331
rect 909 331 915 347
rect 931 359 935 436
rect 1005 359 1009 436
rect 931 347 934 359
rect 1006 347 1009 359
rect 931 331 937 347
rect 909 324 917 331
rect 863 304 867 324
rect 913 304 917 324
rect 923 324 937 331
rect 1003 331 1009 347
rect 1025 359 1029 436
rect 1085 359 1089 436
rect 1025 347 1034 359
rect 1086 347 1089 359
rect 1025 331 1031 347
rect 1003 324 1017 331
rect 923 304 927 324
rect 1013 304 1017 324
rect 1023 324 1031 331
rect 1083 331 1089 347
rect 1105 359 1109 436
rect 1165 373 1169 396
rect 1166 361 1169 373
rect 1105 347 1114 359
rect 1105 331 1111 347
rect 1083 324 1097 331
rect 1023 304 1027 324
rect 1093 304 1097 324
rect 1103 324 1111 331
rect 1103 304 1107 324
rect 1160 313 1166 361
rect 1185 339 1189 396
rect 1205 374 1209 396
rect 1225 374 1229 396
rect 1276 392 1280 396
rect 1262 384 1280 392
rect 1205 368 1218 374
rect 1225 373 1245 374
rect 1262 373 1266 384
rect 1225 368 1233 373
rect 1214 339 1218 368
rect 1187 327 1189 339
rect 1185 325 1189 327
rect 1185 318 1198 325
rect 1160 309 1190 313
rect 1186 304 1190 309
rect 1194 304 1198 318
rect 1214 304 1218 327
rect 1233 319 1239 361
rect 1222 312 1239 319
rect 1262 316 1266 361
rect 1284 339 1288 396
rect 1306 393 1310 436
rect 1306 381 1313 393
rect 1286 327 1295 339
rect 1222 304 1226 312
rect 1262 309 1275 316
rect 1271 304 1275 309
rect 1291 304 1295 327
rect 1311 304 1315 381
rect 1397 373 1401 396
rect 1386 361 1401 373
rect 1405 373 1409 396
rect 1456 392 1460 396
rect 1442 384 1460 392
rect 1442 373 1446 384
rect 1405 361 1414 373
rect 1385 284 1389 361
rect 1405 284 1409 361
rect 1442 316 1446 361
rect 1464 339 1468 396
rect 1486 393 1490 436
rect 1486 381 1493 393
rect 1466 327 1475 339
rect 1442 309 1455 316
rect 1451 304 1455 309
rect 1471 304 1475 327
rect 1491 304 1495 381
rect 1551 353 1555 436
rect 1546 341 1555 353
rect 1551 284 1555 341
rect 1625 339 1629 396
rect 1645 382 1649 396
rect 1665 382 1669 396
rect 1645 376 1660 382
rect 1665 376 1681 382
rect 1654 353 1660 376
rect 1625 327 1634 339
rect 1632 284 1636 327
rect 1654 304 1658 341
rect 1674 339 1681 376
rect 1711 353 1715 436
rect 1771 428 1775 436
rect 1760 424 1775 428
rect 1791 424 1795 436
rect 1760 393 1766 424
rect 1780 420 1795 424
rect 1780 413 1786 420
rect 1766 381 1776 393
rect 1706 341 1715 353
rect 1674 314 1681 327
rect 1662 308 1681 314
rect 1662 304 1666 308
rect 1711 284 1715 341
rect 1772 324 1776 381
rect 1780 324 1784 401
rect 1811 393 1815 436
rect 1788 381 1795 393
rect 1807 381 1815 393
rect 1871 382 1875 396
rect 1891 382 1895 396
rect 1788 324 1792 381
rect 1859 376 1875 382
rect 1880 376 1895 382
rect 1859 339 1866 376
rect 1880 353 1886 376
rect 1859 314 1866 327
rect 1859 308 1878 314
rect 1874 304 1878 308
rect 1882 304 1886 341
rect 1911 339 1915 396
rect 1971 359 1975 436
rect 1966 347 1975 359
rect 1906 327 1915 339
rect 1969 331 1975 347
rect 1991 359 1995 436
rect 2051 359 2055 436
rect 1991 347 1994 359
rect 2046 347 2055 359
rect 1991 331 1997 347
rect 1904 284 1908 327
rect 1969 324 1977 331
rect 1973 304 1977 324
rect 1983 324 1997 331
rect 2049 331 2055 347
rect 2071 359 2075 436
rect 2131 359 2135 436
rect 2071 347 2074 359
rect 2126 347 2135 359
rect 2071 331 2077 347
rect 2049 324 2057 331
rect 1983 304 1987 324
rect 2053 304 2057 324
rect 2063 324 2077 331
rect 2129 331 2135 347
rect 2151 359 2155 436
rect 2237 373 2241 396
rect 2226 361 2241 373
rect 2245 373 2249 396
rect 2245 361 2254 373
rect 2151 347 2154 359
rect 2151 331 2157 347
rect 2129 324 2137 331
rect 2063 304 2067 324
rect 2133 304 2137 324
rect 2143 324 2157 331
rect 2143 304 2147 324
rect 2225 284 2229 361
rect 2245 284 2249 361
rect 2305 359 2309 436
rect 2306 347 2309 359
rect 2303 331 2309 347
rect 2325 359 2329 436
rect 2451 428 2455 436
rect 2440 424 2455 428
rect 2471 424 2475 436
rect 2371 373 2375 396
rect 2366 361 2375 373
rect 2379 373 2383 396
rect 2440 393 2446 424
rect 2460 420 2475 424
rect 2460 413 2466 420
rect 2446 381 2456 393
rect 2379 361 2394 373
rect 2325 347 2334 359
rect 2325 331 2331 347
rect 2303 324 2317 331
rect 2313 304 2317 324
rect 2323 324 2331 331
rect 2323 304 2327 324
rect 2371 284 2375 361
rect 2391 284 2395 361
rect 2452 324 2456 381
rect 2460 324 2464 401
rect 2491 393 2495 436
rect 2468 381 2475 393
rect 2487 381 2495 393
rect 2468 324 2472 381
rect 2565 353 2569 436
rect 2625 393 2629 436
rect 2645 424 2649 436
rect 2665 428 2669 436
rect 2665 424 2680 428
rect 2645 420 2660 424
rect 2654 413 2660 420
rect 2625 381 2633 393
rect 2645 381 2652 393
rect 2565 341 2574 353
rect 2565 284 2569 341
rect 2648 324 2652 381
rect 2656 324 2660 401
rect 2674 393 2680 424
rect 2664 381 2674 393
rect 2711 382 2715 396
rect 2731 382 2735 396
rect 2664 324 2668 381
rect 2699 376 2715 382
rect 2720 376 2735 382
rect 2699 339 2706 376
rect 2720 353 2726 376
rect 2699 314 2706 327
rect 2699 308 2718 314
rect 2714 304 2718 308
rect 2722 304 2726 341
rect 2751 339 2755 396
rect 2811 373 2815 396
rect 2806 361 2815 373
rect 2819 373 2823 396
rect 2819 361 2834 373
rect 2746 327 2755 339
rect 2744 284 2748 327
rect 2811 284 2815 361
rect 2831 284 2835 361
rect 2905 359 2909 436
rect 2906 347 2909 359
rect 2903 331 2909 347
rect 2925 359 2929 436
rect 2990 393 2994 436
rect 2987 381 2994 393
rect 2925 347 2934 359
rect 2925 331 2931 347
rect 2903 324 2917 331
rect 2913 304 2917 324
rect 2923 324 2931 331
rect 2923 304 2927 324
rect 2985 304 2989 381
rect 3012 339 3016 396
rect 3020 392 3024 396
rect 3090 393 3094 436
rect 3020 384 3038 392
rect 3034 373 3038 384
rect 3087 381 3094 393
rect 3005 327 3014 339
rect 3005 304 3009 327
rect 3034 316 3038 361
rect 3025 309 3038 316
rect 3025 304 3029 309
rect 3085 304 3089 381
rect 3112 339 3116 396
rect 3120 392 3124 396
rect 3120 384 3138 392
rect 3134 373 3138 384
rect 3197 373 3201 396
rect 3186 361 3201 373
rect 3205 373 3209 396
rect 3205 361 3214 373
rect 3105 327 3114 339
rect 3105 304 3109 327
rect 3134 316 3138 361
rect 3125 309 3138 316
rect 3125 304 3129 309
rect 3185 284 3189 361
rect 3205 284 3209 361
rect 3265 353 3269 436
rect 3330 393 3334 436
rect 3327 381 3334 393
rect 3265 341 3274 353
rect 3265 284 3269 341
rect 3325 304 3329 381
rect 3352 339 3356 396
rect 3360 392 3364 396
rect 3360 384 3378 392
rect 3374 373 3378 384
rect 3345 327 3354 339
rect 3345 304 3349 327
rect 3374 316 3378 361
rect 3425 339 3429 396
rect 3445 382 3449 396
rect 3465 382 3469 396
rect 3445 376 3460 382
rect 3465 376 3481 382
rect 3454 353 3460 376
rect 3425 327 3434 339
rect 3365 309 3378 316
rect 3365 304 3369 309
rect 3432 284 3436 327
rect 3454 304 3458 341
rect 3474 339 3481 376
rect 3537 373 3541 396
rect 3526 361 3541 373
rect 3545 373 3549 396
rect 3591 392 3595 396
rect 3582 387 3595 392
rect 3545 361 3554 373
rect 3474 314 3481 327
rect 3462 308 3481 314
rect 3462 304 3466 308
rect 3525 284 3529 361
rect 3545 284 3549 361
rect 3582 353 3586 387
rect 3601 373 3605 396
rect 3621 391 3625 396
rect 3582 296 3586 341
rect 3601 297 3605 361
rect 3691 359 3695 436
rect 3686 347 3695 359
rect 3689 331 3695 347
rect 3711 359 3715 436
rect 3771 359 3775 436
rect 3711 347 3714 359
rect 3766 347 3775 359
rect 3711 331 3717 347
rect 3689 324 3697 331
rect 3625 312 3635 324
rect 3631 304 3635 312
rect 3693 304 3697 324
rect 3703 324 3717 331
rect 3769 331 3775 347
rect 3791 359 3795 436
rect 3870 393 3874 436
rect 3867 381 3874 393
rect 3791 347 3794 359
rect 3791 331 3797 347
rect 3769 324 3777 331
rect 3703 304 3707 324
rect 3773 304 3777 324
rect 3783 324 3797 331
rect 3783 304 3787 324
rect 3865 304 3869 381
rect 3892 339 3896 396
rect 3900 392 3904 396
rect 3900 384 3918 392
rect 3914 373 3918 384
rect 3885 327 3894 339
rect 3885 304 3889 327
rect 3914 316 3918 361
rect 3905 309 3918 316
rect 3965 353 3969 436
rect 4025 353 4029 436
rect 4093 433 4097 456
rect 4089 426 4097 433
rect 4089 397 4093 426
rect 4101 416 4105 456
rect 4121 404 4125 436
rect 4129 432 4133 436
rect 4129 430 4165 432
rect 4129 428 4153 430
rect 4071 384 4075 396
rect 4089 391 4097 397
rect 4071 372 4073 384
rect 3965 341 3974 353
rect 4025 341 4034 353
rect 3905 304 3909 309
rect 3582 291 3595 296
rect 3601 291 3615 297
rect 3591 284 3595 291
rect 3611 284 3615 291
rect 3965 284 3969 341
rect 4025 284 4029 341
rect 4071 304 4075 372
rect 4093 345 4097 391
rect 4093 284 4097 333
rect 4121 309 4127 404
rect 4103 305 4127 309
rect 4103 284 4107 305
rect 4123 300 4141 301
rect 4123 296 4153 300
rect 4123 284 4127 296
rect 4161 292 4165 418
rect 4175 410 4179 436
rect 4195 430 4199 436
rect 4131 288 4165 292
rect 4131 284 4135 288
rect 4177 284 4181 398
rect 4193 308 4197 418
rect 4207 396 4211 436
rect 4202 384 4205 396
rect 4202 320 4206 384
rect 4227 377 4231 436
rect 4222 369 4231 377
rect 4222 340 4226 369
rect 4241 354 4245 436
rect 4261 353 4265 396
rect 4325 359 4329 436
rect 4202 316 4235 320
rect 4201 296 4203 308
rect 4199 284 4203 296
rect 4209 296 4211 308
rect 4209 284 4213 296
rect 4231 284 4235 316
rect 4241 284 4245 342
rect 4326 347 4329 359
rect 4261 304 4265 341
rect 4323 331 4329 347
rect 4345 359 4349 436
rect 4410 393 4414 436
rect 4407 381 4414 393
rect 4345 347 4354 359
rect 4345 331 4351 347
rect 4323 324 4337 331
rect 4333 304 4337 324
rect 4343 324 4351 331
rect 4343 304 4347 324
rect 4405 304 4409 381
rect 4432 339 4436 396
rect 4440 392 4444 396
rect 4440 384 4458 392
rect 4454 373 4458 384
rect 4425 327 4434 339
rect 4425 304 4429 327
rect 4454 316 4458 361
rect 4445 309 4458 316
rect 4505 353 4509 436
rect 4573 433 4577 456
rect 4569 426 4577 433
rect 4569 397 4573 426
rect 4581 416 4585 456
rect 4601 404 4605 436
rect 4609 432 4613 436
rect 4609 430 4645 432
rect 4609 428 4633 430
rect 4551 384 4555 396
rect 4569 391 4577 397
rect 4551 372 4553 384
rect 4505 341 4514 353
rect 4445 304 4449 309
rect 4505 284 4509 341
rect 4551 304 4555 372
rect 4573 345 4577 391
rect 4573 284 4577 333
rect 4601 309 4607 404
rect 4583 305 4607 309
rect 4583 284 4587 305
rect 4603 300 4621 301
rect 4603 296 4633 300
rect 4603 284 4607 296
rect 4641 292 4645 418
rect 4655 410 4659 436
rect 4675 430 4679 436
rect 4611 288 4645 292
rect 4611 284 4615 288
rect 4657 284 4661 398
rect 4673 308 4677 418
rect 4687 396 4691 436
rect 4682 384 4685 396
rect 4682 320 4686 384
rect 4707 377 4711 436
rect 4702 369 4711 377
rect 4702 340 4706 369
rect 4721 354 4725 436
rect 4741 353 4745 396
rect 4682 316 4715 320
rect 4681 296 4683 308
rect 4679 284 4683 296
rect 4689 296 4691 308
rect 4689 284 4693 296
rect 4711 284 4715 316
rect 4721 284 4725 342
rect 4741 304 4745 341
rect 33 260 37 264
rect 43 260 47 264
rect 113 260 117 264
rect 123 260 127 264
rect 213 260 217 264
rect 223 260 227 264
rect 293 260 297 264
rect 303 260 307 264
rect 375 260 379 264
rect 395 260 399 264
rect 405 260 409 264
rect 473 260 477 264
rect 483 260 487 264
rect 568 260 572 264
rect 576 260 580 264
rect 584 260 588 264
rect 666 260 670 264
rect 674 260 678 264
rect 694 260 698 264
rect 702 260 706 264
rect 765 260 769 264
rect 785 260 789 264
rect 853 260 857 264
rect 863 260 867 264
rect 913 260 917 264
rect 923 260 927 264
rect 1013 260 1017 264
rect 1023 260 1027 264
rect 1093 260 1097 264
rect 1103 260 1107 264
rect 1186 260 1190 264
rect 1194 260 1198 264
rect 1214 260 1218 264
rect 1222 260 1226 264
rect 1271 260 1275 264
rect 1291 260 1295 264
rect 1311 260 1315 264
rect 1385 260 1389 264
rect 1405 260 1409 264
rect 1451 260 1455 264
rect 1471 260 1475 264
rect 1491 260 1495 264
rect 1551 260 1555 264
rect 1632 260 1636 264
rect 1654 260 1658 264
rect 1662 260 1666 264
rect 1711 260 1715 264
rect 1772 260 1776 264
rect 1780 260 1784 264
rect 1788 260 1792 264
rect 1874 260 1878 264
rect 1882 260 1886 264
rect 1904 260 1908 264
rect 1973 260 1977 264
rect 1983 260 1987 264
rect 2053 260 2057 264
rect 2063 260 2067 264
rect 2133 260 2137 264
rect 2143 260 2147 264
rect 2225 260 2229 264
rect 2245 260 2249 264
rect 2313 260 2317 264
rect 2323 260 2327 264
rect 2371 260 2375 264
rect 2391 260 2395 264
rect 2452 260 2456 264
rect 2460 260 2464 264
rect 2468 260 2472 264
rect 2565 260 2569 264
rect 2648 260 2652 264
rect 2656 260 2660 264
rect 2664 260 2668 264
rect 2714 260 2718 264
rect 2722 260 2726 264
rect 2744 260 2748 264
rect 2811 260 2815 264
rect 2831 260 2835 264
rect 2913 260 2917 264
rect 2923 260 2927 264
rect 2985 260 2989 264
rect 3005 260 3009 264
rect 3025 260 3029 264
rect 3085 260 3089 264
rect 3105 260 3109 264
rect 3125 260 3129 264
rect 3185 260 3189 264
rect 3205 260 3209 264
rect 3265 260 3269 264
rect 3325 260 3329 264
rect 3345 260 3349 264
rect 3365 260 3369 264
rect 3432 260 3436 264
rect 3454 260 3458 264
rect 3462 260 3466 264
rect 3525 260 3529 264
rect 3545 260 3549 264
rect 3591 260 3595 264
rect 3611 260 3615 264
rect 3631 260 3635 264
rect 3693 260 3697 264
rect 3703 260 3707 264
rect 3773 260 3777 264
rect 3783 260 3787 264
rect 3865 260 3869 264
rect 3885 260 3889 264
rect 3905 260 3909 264
rect 3965 260 3969 264
rect 4025 260 4029 264
rect 4071 260 4075 264
rect 4093 260 4097 264
rect 4103 260 4107 264
rect 4123 260 4127 264
rect 4131 260 4135 264
rect 4177 260 4181 264
rect 4199 260 4203 264
rect 4209 260 4213 264
rect 4231 260 4235 264
rect 4241 260 4245 264
rect 4261 260 4265 264
rect 4333 260 4337 264
rect 4343 260 4347 264
rect 4405 260 4409 264
rect 4425 260 4429 264
rect 4445 260 4449 264
rect 4505 260 4509 264
rect 4551 260 4555 264
rect 4573 260 4577 264
rect 4583 260 4587 264
rect 4603 260 4607 264
rect 4611 260 4615 264
rect 4657 260 4661 264
rect 4679 260 4683 264
rect 4689 260 4693 264
rect 4711 260 4715 264
rect 4721 260 4725 264
rect 4741 260 4745 264
rect 68 236 72 240
rect 76 236 80 240
rect 84 236 88 240
rect 134 236 138 240
rect 142 236 146 240
rect 164 236 168 240
rect 245 236 249 240
rect 265 236 269 240
rect 285 236 289 240
rect 331 236 335 240
rect 351 236 355 240
rect 371 236 375 240
rect 468 236 472 240
rect 476 236 480 240
rect 484 236 488 240
rect 532 236 536 240
rect 540 236 544 240
rect 548 236 552 240
rect 634 236 638 240
rect 642 236 646 240
rect 664 236 668 240
rect 752 236 756 240
rect 774 236 778 240
rect 782 236 786 240
rect 831 236 835 240
rect 905 236 909 240
rect 925 236 929 240
rect 945 236 949 240
rect 1005 236 1009 240
rect 1051 236 1055 240
rect 1071 236 1075 240
rect 1091 236 1095 240
rect 1151 236 1155 240
rect 1171 236 1175 240
rect 1191 236 1195 240
rect 1252 236 1256 240
rect 1260 236 1264 240
rect 1268 236 1272 240
rect 1352 236 1356 240
rect 1360 236 1364 240
rect 1368 236 1372 240
rect 1472 236 1476 240
rect 1494 236 1498 240
rect 1502 236 1506 240
rect 1552 236 1556 240
rect 1560 236 1564 240
rect 1568 236 1572 240
rect 1672 236 1676 240
rect 1694 236 1698 240
rect 1702 236 1706 240
rect 1752 236 1756 240
rect 1760 236 1764 240
rect 1768 236 1772 240
rect 1853 236 1857 240
rect 1863 236 1867 240
rect 1931 236 1935 240
rect 1953 236 1957 240
rect 2035 236 2039 240
rect 2055 236 2059 240
rect 2065 236 2069 240
rect 2111 236 2115 240
rect 2133 236 2137 240
rect 2192 236 2196 240
rect 2200 236 2204 240
rect 2208 236 2212 240
rect 2294 236 2298 240
rect 2302 236 2306 240
rect 2322 236 2326 240
rect 2330 236 2334 240
rect 2411 236 2415 240
rect 2431 236 2435 240
rect 2451 236 2455 240
rect 2532 236 2536 240
rect 2554 236 2558 240
rect 2562 236 2566 240
rect 2611 236 2615 240
rect 2631 236 2635 240
rect 2651 236 2655 240
rect 2711 236 2715 240
rect 2772 236 2776 240
rect 2780 236 2784 240
rect 2788 236 2792 240
rect 2871 236 2875 240
rect 2935 236 2939 240
rect 2955 236 2959 240
rect 2965 236 2969 240
rect 2987 236 2991 240
rect 2997 236 3001 240
rect 3019 236 3023 240
rect 3065 236 3069 240
rect 3073 236 3077 240
rect 3093 236 3097 240
rect 3103 236 3107 240
rect 3125 236 3129 240
rect 3171 236 3175 240
rect 3245 236 3249 240
rect 3295 236 3299 240
rect 3315 236 3319 240
rect 3325 236 3329 240
rect 3347 236 3351 240
rect 3357 236 3361 240
rect 3379 236 3383 240
rect 3425 236 3429 240
rect 3433 236 3437 240
rect 3453 236 3457 240
rect 3463 236 3467 240
rect 3485 236 3489 240
rect 3545 236 3549 240
rect 3565 236 3569 240
rect 3611 236 3615 240
rect 3633 236 3637 240
rect 3643 236 3647 240
rect 3663 236 3667 240
rect 3671 236 3675 240
rect 3717 236 3721 240
rect 3739 236 3743 240
rect 3749 236 3753 240
rect 3771 236 3775 240
rect 3781 236 3785 240
rect 3801 236 3805 240
rect 3851 236 3855 240
rect 3911 236 3915 240
rect 3931 236 3935 240
rect 3951 236 3955 240
rect 4011 236 4015 240
rect 4031 236 4035 240
rect 4091 236 4095 240
rect 4111 236 4115 240
rect 4185 236 4189 240
rect 4205 236 4209 240
rect 4251 236 4255 240
rect 4271 236 4275 240
rect 4291 236 4295 240
rect 4373 236 4377 240
rect 4383 236 4387 240
rect 4445 236 4449 240
rect 4491 236 4495 240
rect 4511 236 4515 240
rect 4573 236 4577 240
rect 4583 236 4587 240
rect 4665 236 4669 240
rect 4713 236 4717 240
rect 4723 236 4727 240
rect 134 192 138 196
rect 119 186 138 192
rect 68 119 72 176
rect 45 107 53 119
rect 65 107 72 119
rect 45 64 49 107
rect 76 99 80 176
rect 84 119 88 176
rect 119 173 126 186
rect 119 124 126 161
rect 142 159 146 196
rect 164 173 168 216
rect 166 161 175 173
rect 140 124 146 147
rect 84 107 94 119
rect 119 118 135 124
rect 140 118 155 124
rect 74 80 80 87
rect 65 76 80 80
rect 94 76 100 107
rect 131 104 135 118
rect 151 104 155 118
rect 171 104 175 161
rect 245 119 249 196
rect 265 173 269 196
rect 285 191 289 196
rect 331 191 335 196
rect 285 184 298 191
rect 265 161 274 173
rect 247 107 254 119
rect 65 64 69 76
rect 85 72 100 76
rect 85 64 89 72
rect 250 64 254 107
rect 272 104 276 161
rect 294 139 298 184
rect 322 184 335 191
rect 322 139 326 184
rect 351 173 355 196
rect 346 161 355 173
rect 294 116 298 127
rect 280 108 298 116
rect 322 116 326 127
rect 322 108 340 116
rect 280 104 284 108
rect 336 104 340 108
rect 344 104 348 161
rect 371 119 375 196
rect 634 192 638 196
rect 619 186 638 192
rect 468 119 472 176
rect 366 107 373 119
rect 445 107 453 119
rect 465 107 472 119
rect 366 64 370 107
rect 445 64 449 107
rect 476 99 480 176
rect 484 119 488 176
rect 532 119 536 176
rect 484 107 494 119
rect 526 107 536 119
rect 474 80 480 87
rect 465 76 480 80
rect 494 76 500 107
rect 465 64 469 76
rect 485 72 500 76
rect 520 76 526 107
rect 540 99 544 176
rect 548 119 552 176
rect 619 173 626 186
rect 619 124 626 161
rect 642 159 646 196
rect 664 173 668 216
rect 752 173 756 216
rect 666 161 675 173
rect 640 124 646 147
rect 548 107 555 119
rect 567 107 575 119
rect 619 118 635 124
rect 640 118 655 124
rect 540 80 546 87
rect 540 76 555 80
rect 520 72 535 76
rect 485 64 489 72
rect 531 64 535 72
rect 551 64 555 76
rect 571 64 575 107
rect 631 104 635 118
rect 651 104 655 118
rect 671 104 675 161
rect 745 161 754 173
rect 745 104 749 161
rect 774 159 778 196
rect 782 192 786 196
rect 782 186 801 192
rect 794 173 801 186
rect 774 124 780 147
rect 794 124 801 161
rect 831 159 835 216
rect 826 147 835 159
rect 765 118 780 124
rect 785 118 801 124
rect 765 104 769 118
rect 785 104 789 118
rect 831 64 835 147
rect 905 119 909 196
rect 925 173 929 196
rect 945 191 949 196
rect 945 184 958 191
rect 925 161 934 173
rect 907 107 914 119
rect 910 64 914 107
rect 932 104 936 161
rect 954 139 958 184
rect 1005 159 1009 216
rect 1051 191 1055 196
rect 1042 184 1055 191
rect 1005 147 1014 159
rect 954 116 958 127
rect 940 108 958 116
rect 940 104 944 108
rect 1005 64 1009 147
rect 1042 139 1046 184
rect 1071 173 1075 196
rect 1066 161 1075 173
rect 1042 116 1046 127
rect 1042 108 1060 116
rect 1056 104 1060 108
rect 1064 104 1068 161
rect 1091 119 1095 196
rect 1151 191 1155 196
rect 1142 184 1155 191
rect 1142 139 1146 184
rect 1171 173 1175 196
rect 1166 161 1175 173
rect 1086 107 1093 119
rect 1142 116 1146 127
rect 1142 108 1160 116
rect 1086 64 1090 107
rect 1156 104 1160 108
rect 1164 104 1168 161
rect 1191 119 1195 196
rect 1252 119 1256 176
rect 1186 107 1193 119
rect 1246 107 1256 119
rect 1186 64 1190 107
rect 1240 76 1246 107
rect 1260 99 1264 176
rect 1268 119 1272 176
rect 1352 119 1356 176
rect 1268 107 1275 119
rect 1287 107 1295 119
rect 1346 107 1356 119
rect 1260 80 1266 87
rect 1260 76 1275 80
rect 1240 72 1255 76
rect 1251 64 1255 72
rect 1271 64 1275 76
rect 1291 64 1295 107
rect 1340 76 1346 107
rect 1360 99 1364 176
rect 1368 119 1372 176
rect 1472 173 1476 216
rect 1465 161 1474 173
rect 1368 107 1375 119
rect 1387 107 1395 119
rect 1360 80 1366 87
rect 1360 76 1375 80
rect 1340 72 1355 76
rect 1351 64 1355 72
rect 1371 64 1375 76
rect 1391 64 1395 107
rect 1465 104 1469 161
rect 1494 159 1498 196
rect 1502 192 1506 196
rect 1502 186 1521 192
rect 1514 173 1521 186
rect 1494 124 1500 147
rect 1514 124 1521 161
rect 1485 118 1500 124
rect 1505 118 1521 124
rect 1552 119 1556 176
rect 1485 104 1489 118
rect 1505 104 1509 118
rect 1546 107 1556 119
rect 1540 76 1546 107
rect 1560 99 1564 176
rect 1568 119 1572 176
rect 1672 173 1676 216
rect 1665 161 1674 173
rect 1568 107 1575 119
rect 1587 107 1595 119
rect 1560 80 1566 87
rect 1560 76 1575 80
rect 1540 72 1555 76
rect 1551 64 1555 72
rect 1571 64 1575 76
rect 1591 64 1595 107
rect 1665 104 1669 161
rect 1694 159 1698 196
rect 1702 192 1706 196
rect 1702 186 1721 192
rect 1714 173 1721 186
rect 1853 176 1857 196
rect 1694 124 1700 147
rect 1714 124 1721 161
rect 1685 118 1700 124
rect 1705 118 1721 124
rect 1752 119 1756 176
rect 1685 104 1689 118
rect 1705 104 1709 118
rect 1746 107 1756 119
rect 1740 76 1746 107
rect 1760 99 1764 176
rect 1768 119 1772 176
rect 1849 169 1857 176
rect 1863 176 1867 196
rect 1863 169 1877 176
rect 1849 153 1855 169
rect 1846 141 1855 153
rect 1768 107 1775 119
rect 1787 107 1795 119
rect 1760 80 1766 87
rect 1760 76 1775 80
rect 1740 72 1755 76
rect 1751 64 1755 72
rect 1771 64 1775 76
rect 1791 64 1795 107
rect 1851 64 1855 141
rect 1871 153 1877 169
rect 1871 141 1874 153
rect 1871 64 1875 141
rect 1931 139 1935 216
rect 1953 190 1957 196
rect 2035 190 2039 196
rect 1955 178 1957 190
rect 2021 178 2033 190
rect 1926 127 1935 139
rect 1931 64 1935 127
rect 1955 110 1957 122
rect 1953 104 1957 110
rect 2021 104 2025 178
rect 2055 153 2059 196
rect 2046 141 2059 153
rect 2043 64 2047 141
rect 2065 139 2069 196
rect 2111 139 2115 216
rect 2133 190 2137 196
rect 2135 178 2137 190
rect 2294 188 2298 196
rect 2281 181 2298 188
rect 2065 127 2074 139
rect 2106 127 2115 139
rect 2065 64 2069 127
rect 2111 64 2115 127
rect 2135 110 2137 122
rect 2192 119 2196 176
rect 2133 104 2137 110
rect 2186 107 2196 119
rect 2180 76 2186 107
rect 2200 99 2204 176
rect 2208 119 2212 176
rect 2281 139 2287 181
rect 2302 173 2306 196
rect 2322 182 2326 196
rect 2330 191 2334 196
rect 2411 191 2415 196
rect 2330 187 2360 191
rect 2322 175 2335 182
rect 2331 173 2335 175
rect 2331 161 2333 173
rect 2302 132 2306 161
rect 2287 127 2295 132
rect 2275 126 2295 127
rect 2302 126 2315 132
rect 2208 107 2215 119
rect 2227 107 2235 119
rect 2200 80 2206 87
rect 2200 76 2215 80
rect 2180 72 2195 76
rect 2191 64 2195 72
rect 2211 64 2215 76
rect 2231 64 2235 107
rect 2291 104 2295 126
rect 2311 104 2315 126
rect 2331 104 2335 161
rect 2354 139 2360 187
rect 2402 184 2415 191
rect 2402 139 2406 184
rect 2431 173 2435 196
rect 2426 161 2435 173
rect 2351 127 2354 139
rect 2351 104 2355 127
rect 2402 116 2406 127
rect 2402 108 2420 116
rect 2416 104 2420 108
rect 2424 104 2428 161
rect 2451 119 2455 196
rect 2532 173 2536 216
rect 2525 161 2534 173
rect 2446 107 2453 119
rect 2446 64 2450 107
rect 2525 104 2529 161
rect 2554 159 2558 196
rect 2562 192 2566 196
rect 2562 186 2581 192
rect 2611 191 2615 196
rect 2574 173 2581 186
rect 2602 184 2615 191
rect 2554 124 2560 147
rect 2574 124 2581 161
rect 2602 139 2606 184
rect 2631 173 2635 196
rect 2626 161 2635 173
rect 2545 118 2560 124
rect 2565 118 2581 124
rect 2545 104 2549 118
rect 2565 104 2569 118
rect 2602 116 2606 127
rect 2602 108 2620 116
rect 2616 104 2620 108
rect 2624 104 2628 161
rect 2651 119 2655 196
rect 2711 159 2715 216
rect 2706 147 2715 159
rect 2646 107 2653 119
rect 2646 64 2650 107
rect 2711 64 2715 147
rect 2772 119 2776 176
rect 2766 107 2776 119
rect 2760 76 2766 107
rect 2780 99 2784 176
rect 2788 119 2792 176
rect 2871 159 2875 216
rect 2935 159 2939 196
rect 2866 147 2875 159
rect 2955 158 2959 216
rect 2965 184 2969 216
rect 2987 204 2991 216
rect 2989 192 2991 204
rect 2997 204 3001 216
rect 2997 192 2999 204
rect 2965 180 2998 184
rect 2788 107 2795 119
rect 2807 107 2815 119
rect 2780 80 2786 87
rect 2780 76 2795 80
rect 2760 72 2775 76
rect 2771 64 2775 72
rect 2791 64 2795 76
rect 2811 64 2815 107
rect 2871 64 2875 147
rect 2935 104 2939 147
rect 2955 64 2959 146
rect 2974 131 2978 160
rect 2969 123 2978 131
rect 2969 64 2973 123
rect 2994 116 2998 180
rect 2995 104 2998 116
rect 2989 64 2993 104
rect 3003 82 3007 192
rect 3019 102 3023 216
rect 3065 212 3069 216
rect 3035 208 3069 212
rect 3001 64 3005 70
rect 3021 64 3025 90
rect 3035 82 3039 208
rect 3073 204 3077 216
rect 3047 200 3077 204
rect 3059 199 3077 200
rect 3093 195 3097 216
rect 3073 191 3097 195
rect 3073 96 3079 191
rect 3103 167 3107 216
rect 3103 109 3107 155
rect 3125 128 3129 196
rect 3171 159 3175 216
rect 3166 147 3175 159
rect 3127 116 3129 128
rect 3103 103 3111 109
rect 3125 104 3129 116
rect 3047 70 3071 72
rect 3035 68 3071 70
rect 3067 64 3071 68
rect 3075 64 3079 96
rect 3095 44 3099 84
rect 3107 74 3111 103
rect 3103 67 3111 74
rect 3103 44 3107 67
rect 3171 64 3175 147
rect 3245 159 3249 216
rect 3295 159 3299 196
rect 3245 147 3254 159
rect 3315 158 3319 216
rect 3325 184 3329 216
rect 3347 204 3351 216
rect 3349 192 3351 204
rect 3357 204 3361 216
rect 3357 192 3359 204
rect 3325 180 3358 184
rect 3245 64 3249 147
rect 3295 104 3299 147
rect 3315 64 3319 146
rect 3334 131 3338 160
rect 3329 123 3338 131
rect 3329 64 3333 123
rect 3354 116 3358 180
rect 3355 104 3358 116
rect 3349 64 3353 104
rect 3363 82 3367 192
rect 3379 102 3383 216
rect 3425 212 3429 216
rect 3395 208 3429 212
rect 3361 64 3365 70
rect 3381 64 3385 90
rect 3395 82 3399 208
rect 3433 204 3437 216
rect 3407 200 3437 204
rect 3419 199 3437 200
rect 3453 195 3457 216
rect 3433 191 3457 195
rect 3433 96 3439 191
rect 3463 167 3467 216
rect 3463 109 3467 155
rect 3485 128 3489 196
rect 3545 139 3549 216
rect 3565 139 3569 216
rect 3487 116 3489 128
rect 3546 127 3561 139
rect 3463 103 3471 109
rect 3485 104 3489 116
rect 3557 104 3561 127
rect 3565 127 3574 139
rect 3611 128 3615 196
rect 3633 167 3637 216
rect 3643 195 3647 216
rect 3663 204 3667 216
rect 3671 212 3675 216
rect 3671 208 3705 212
rect 3663 200 3693 204
rect 3663 199 3681 200
rect 3643 191 3667 195
rect 3565 104 3569 127
rect 3611 116 3613 128
rect 3611 104 3615 116
rect 3633 109 3637 155
rect 3407 70 3431 72
rect 3395 68 3431 70
rect 3427 64 3431 68
rect 3435 64 3439 96
rect 3455 44 3459 84
rect 3467 74 3471 103
rect 3463 67 3471 74
rect 3463 44 3467 67
rect 3629 103 3637 109
rect 3629 74 3633 103
rect 3661 96 3667 191
rect 3629 67 3637 74
rect 3633 44 3637 67
rect 3641 44 3645 84
rect 3661 64 3665 96
rect 3701 82 3705 208
rect 3717 102 3721 216
rect 3739 204 3743 216
rect 3741 192 3743 204
rect 3749 204 3753 216
rect 3749 192 3751 204
rect 3669 70 3693 72
rect 3669 68 3705 70
rect 3669 64 3673 68
rect 3715 64 3719 90
rect 3733 82 3737 192
rect 3771 184 3775 216
rect 3742 180 3775 184
rect 3742 116 3746 180
rect 3762 131 3766 160
rect 3781 158 3785 216
rect 3801 159 3805 196
rect 3851 159 3855 216
rect 3911 191 3915 196
rect 3846 147 3855 159
rect 3762 123 3771 131
rect 3742 104 3745 116
rect 3735 64 3739 70
rect 3747 64 3751 104
rect 3767 64 3771 123
rect 3781 64 3785 146
rect 3801 104 3805 147
rect 3851 64 3855 147
rect 3902 184 3915 191
rect 3902 139 3906 184
rect 3931 173 3935 196
rect 3926 161 3935 173
rect 3902 116 3906 127
rect 3902 108 3920 116
rect 3916 104 3920 108
rect 3924 104 3928 161
rect 3951 119 3955 196
rect 4011 139 4015 216
rect 4031 139 4035 216
rect 4091 139 4095 216
rect 4111 139 4115 216
rect 4185 139 4189 216
rect 4205 139 4209 216
rect 4251 191 4255 196
rect 4242 184 4255 191
rect 4242 139 4246 184
rect 4271 173 4275 196
rect 4266 161 4275 173
rect 4006 127 4015 139
rect 3946 107 3953 119
rect 3946 64 3950 107
rect 4011 104 4015 127
rect 4019 127 4034 139
rect 4086 127 4095 139
rect 4019 104 4023 127
rect 4091 104 4095 127
rect 4099 127 4114 139
rect 4186 127 4201 139
rect 4099 104 4103 127
rect 4197 104 4201 127
rect 4205 127 4214 139
rect 4205 104 4209 127
rect 4242 116 4246 127
rect 4242 108 4260 116
rect 4256 104 4260 108
rect 4264 104 4268 161
rect 4291 119 4295 196
rect 4373 176 4377 196
rect 4363 169 4377 176
rect 4383 176 4387 196
rect 4383 169 4391 176
rect 4363 153 4369 169
rect 4366 141 4369 153
rect 4286 107 4293 119
rect 4286 64 4290 107
rect 4365 64 4369 141
rect 4385 153 4391 169
rect 4445 159 4449 216
rect 4385 141 4394 153
rect 4445 147 4454 159
rect 4385 64 4389 141
rect 4445 64 4449 147
rect 4491 139 4495 216
rect 4511 139 4515 216
rect 4573 176 4577 196
rect 4569 169 4577 176
rect 4583 176 4587 196
rect 4583 169 4597 176
rect 4569 153 4575 169
rect 4566 141 4575 153
rect 4486 127 4495 139
rect 4491 104 4495 127
rect 4499 127 4514 139
rect 4499 104 4503 127
rect 4571 64 4575 141
rect 4591 153 4597 169
rect 4665 159 4669 216
rect 4713 176 4717 196
rect 4709 169 4717 176
rect 4723 176 4727 196
rect 4723 169 4737 176
rect 4591 141 4594 153
rect 4665 147 4674 159
rect 4709 153 4715 169
rect 4591 64 4595 141
rect 4665 64 4669 147
rect 4706 141 4715 153
rect 4711 64 4715 141
rect 4731 153 4737 169
rect 4731 141 4734 153
rect 4731 64 4735 141
rect 45 20 49 24
rect 65 20 69 24
rect 85 20 89 24
rect 131 20 135 24
rect 151 20 155 24
rect 171 20 175 24
rect 250 20 254 24
rect 272 20 276 24
rect 280 20 284 24
rect 336 20 340 24
rect 344 20 348 24
rect 366 20 370 24
rect 445 20 449 24
rect 465 20 469 24
rect 485 20 489 24
rect 531 20 535 24
rect 551 20 555 24
rect 571 20 575 24
rect 631 20 635 24
rect 651 20 655 24
rect 671 20 675 24
rect 745 20 749 24
rect 765 20 769 24
rect 785 20 789 24
rect 831 20 835 24
rect 910 20 914 24
rect 932 20 936 24
rect 940 20 944 24
rect 1005 20 1009 24
rect 1056 20 1060 24
rect 1064 20 1068 24
rect 1086 20 1090 24
rect 1156 20 1160 24
rect 1164 20 1168 24
rect 1186 20 1190 24
rect 1251 20 1255 24
rect 1271 20 1275 24
rect 1291 20 1295 24
rect 1351 20 1355 24
rect 1371 20 1375 24
rect 1391 20 1395 24
rect 1465 20 1469 24
rect 1485 20 1489 24
rect 1505 20 1509 24
rect 1551 20 1555 24
rect 1571 20 1575 24
rect 1591 20 1595 24
rect 1665 20 1669 24
rect 1685 20 1689 24
rect 1705 20 1709 24
rect 1751 20 1755 24
rect 1771 20 1775 24
rect 1791 20 1795 24
rect 1851 20 1855 24
rect 1871 20 1875 24
rect 1931 20 1935 24
rect 1953 20 1957 24
rect 2021 20 2025 24
rect 2043 20 2047 24
rect 2065 20 2069 24
rect 2111 20 2115 24
rect 2133 20 2137 24
rect 2191 20 2195 24
rect 2211 20 2215 24
rect 2231 20 2235 24
rect 2291 20 2295 24
rect 2311 20 2315 24
rect 2331 20 2335 24
rect 2351 20 2355 24
rect 2416 20 2420 24
rect 2424 20 2428 24
rect 2446 20 2450 24
rect 2525 20 2529 24
rect 2545 20 2549 24
rect 2565 20 2569 24
rect 2616 20 2620 24
rect 2624 20 2628 24
rect 2646 20 2650 24
rect 2711 20 2715 24
rect 2771 20 2775 24
rect 2791 20 2795 24
rect 2811 20 2815 24
rect 2871 20 2875 24
rect 2935 20 2939 24
rect 2955 20 2959 24
rect 2969 20 2973 24
rect 2989 20 2993 24
rect 3001 20 3005 24
rect 3021 20 3025 24
rect 3067 20 3071 24
rect 3075 20 3079 24
rect 3095 20 3099 24
rect 3103 20 3107 24
rect 3125 20 3129 24
rect 3171 20 3175 24
rect 3245 20 3249 24
rect 3295 20 3299 24
rect 3315 20 3319 24
rect 3329 20 3333 24
rect 3349 20 3353 24
rect 3361 20 3365 24
rect 3381 20 3385 24
rect 3427 20 3431 24
rect 3435 20 3439 24
rect 3455 20 3459 24
rect 3463 20 3467 24
rect 3485 20 3489 24
rect 3557 20 3561 24
rect 3565 20 3569 24
rect 3611 20 3615 24
rect 3633 20 3637 24
rect 3641 20 3645 24
rect 3661 20 3665 24
rect 3669 20 3673 24
rect 3715 20 3719 24
rect 3735 20 3739 24
rect 3747 20 3751 24
rect 3767 20 3771 24
rect 3781 20 3785 24
rect 3801 20 3805 24
rect 3851 20 3855 24
rect 3916 20 3920 24
rect 3924 20 3928 24
rect 3946 20 3950 24
rect 4011 20 4015 24
rect 4019 20 4023 24
rect 4091 20 4095 24
rect 4099 20 4103 24
rect 4197 20 4201 24
rect 4205 20 4209 24
rect 4256 20 4260 24
rect 4264 20 4268 24
rect 4286 20 4290 24
rect 4365 20 4369 24
rect 4385 20 4389 24
rect 4445 20 4449 24
rect 4491 20 4495 24
rect 4499 20 4503 24
rect 4571 20 4575 24
rect 4591 20 4595 24
rect 4665 20 4669 24
rect 4711 20 4715 24
rect 4731 20 4735 24
<< polycontact >>
rect 54 4481 66 4493
rect 94 4481 106 4493
rect 74 4467 86 4479
rect 153 4427 165 4439
rect 194 4427 206 4439
rect 214 4427 226 4439
rect 174 4407 186 4419
rect 255 4427 267 4439
rect 234 4407 246 4419
rect 353 4427 365 4439
rect 414 4481 426 4493
rect 454 4481 466 4493
rect 434 4467 446 4479
rect 394 4427 406 4439
rect 374 4407 386 4419
rect 534 4481 546 4493
rect 514 4447 526 4459
rect 634 4481 646 4493
rect 614 4447 626 4459
rect 573 4427 585 4439
rect 673 4427 685 4439
rect 753 4427 765 4439
rect 794 4427 806 4439
rect 814 4427 826 4439
rect 774 4407 786 4419
rect 914 4461 926 4473
rect 855 4427 867 4439
rect 834 4407 846 4419
rect 954 4461 966 4473
rect 994 4427 1006 4439
rect 1094 4481 1106 4493
rect 1134 4481 1146 4493
rect 1114 4467 1126 4479
rect 1035 4427 1047 4439
rect 1014 4407 1026 4419
rect 1214 4461 1226 4473
rect 1254 4461 1266 4473
rect 1294 4447 1306 4459
rect 1334 4447 1346 4459
rect 1414 4481 1426 4493
rect 1375 4427 1387 4439
rect 1474 4461 1486 4473
rect 1434 4447 1446 4459
rect 1514 4461 1526 4473
rect 1534 4447 1546 4459
rect 1574 4447 1586 4459
rect 1614 4427 1626 4439
rect 1754 4481 1766 4493
rect 1655 4427 1667 4439
rect 1634 4407 1646 4419
rect 1794 4481 1806 4493
rect 1774 4467 1786 4479
rect 1814 4467 1826 4479
rect 1934 4481 1946 4493
rect 1914 4467 1926 4479
rect 1974 4481 1986 4493
rect 1954 4467 1966 4479
rect 2114 4467 2126 4479
rect 2034 4447 2046 4459
rect 2074 4447 2086 4459
rect 2194 4481 2206 4493
rect 2174 4447 2186 4459
rect 2318 4481 2330 4493
rect 2354 4481 2366 4493
rect 2295 4447 2307 4459
rect 2233 4427 2245 4439
rect 2394 4467 2406 4479
rect 2374 4447 2386 4459
rect 2433 4496 2445 4508
rect 2494 4481 2506 4493
rect 2414 4447 2426 4459
rect 2534 4481 2546 4493
rect 2514 4467 2526 4479
rect 2433 4429 2445 4441
rect 2635 4481 2647 4493
rect 2673 4481 2685 4493
rect 2614 4447 2626 4459
rect 2734 4467 2746 4479
rect 2777 4512 2789 4524
rect 2799 4512 2811 4524
rect 2774 4480 2786 4492
rect 2693 4447 2705 4459
rect 2754 4466 2766 4478
rect 2783 4424 2795 4436
rect 2815 4410 2827 4422
rect 2801 4390 2813 4402
rect 2847 4508 2859 4520
rect 2901 4475 2913 4487
rect 2915 4436 2927 4448
rect 2994 4467 3006 4479
rect 2863 4404 2875 4416
rect 2835 4390 2847 4402
rect 2887 4404 2899 4416
rect 3074 4481 3086 4493
rect 3035 4427 3047 4439
rect 3094 4447 3106 4459
rect 3134 4447 3146 4459
rect 3174 4447 3186 4459
rect 3254 4481 3266 4493
rect 3215 4427 3227 4439
rect 3414 4467 3426 4479
rect 3274 4447 3286 4459
rect 3314 4447 3326 4459
rect 3354 4447 3366 4459
rect 3467 4475 3479 4487
rect 3453 4436 3465 4448
rect 3521 4508 3533 4520
rect 3481 4404 3493 4416
rect 3505 4404 3517 4416
rect 3569 4512 3581 4524
rect 3591 4512 3603 4524
rect 3553 4410 3565 4422
rect 3533 4390 3545 4402
rect 3594 4480 3606 4492
rect 3614 4466 3626 4478
rect 3634 4467 3646 4479
rect 3585 4424 3597 4436
rect 3567 4390 3579 4402
rect 3694 4481 3706 4493
rect 3674 4447 3686 4459
rect 3774 4461 3786 4473
rect 3733 4427 3745 4439
rect 3898 4484 3910 4496
rect 3938 4484 3950 4496
rect 3978 4484 3990 4496
rect 4085 4498 4097 4510
rect 3814 4461 3826 4473
rect 4014 4481 4026 4493
rect 4134 4461 4146 4473
rect 4114 4447 4126 4459
rect 4085 4430 4097 4442
rect 4174 4461 4186 4473
rect 4214 4467 4226 4479
rect 4294 4481 4306 4493
rect 4274 4447 4286 4459
rect 4407 4475 4419 4487
rect 4333 4427 4345 4439
rect 4393 4436 4405 4448
rect 4461 4508 4473 4520
rect 4421 4404 4433 4416
rect 4445 4404 4457 4416
rect 4509 4512 4521 4524
rect 4531 4512 4543 4524
rect 4493 4410 4505 4422
rect 4473 4390 4485 4402
rect 4534 4480 4546 4492
rect 4554 4466 4566 4478
rect 4574 4467 4586 4479
rect 4525 4424 4537 4436
rect 4507 4390 4519 4402
rect 4643 4498 4655 4510
rect 4694 4461 4706 4473
rect 4614 4447 4626 4459
rect 4643 4430 4655 4442
rect 4734 4461 4746 4473
rect 34 4187 46 4199
rect 74 4187 86 4199
rect 114 4181 126 4193
rect 94 4167 106 4179
rect 214 4187 226 4199
rect 134 4167 146 4179
rect 294 4201 306 4213
rect 375 4221 387 4233
rect 334 4201 346 4213
rect 254 4187 266 4199
rect 434 4201 446 4213
rect 454 4201 466 4213
rect 414 4167 426 4179
rect 513 4221 525 4233
rect 474 4167 486 4179
rect 594 4181 606 4193
rect 674 4181 686 4193
rect 654 4167 666 4179
rect 794 4241 806 4253
rect 774 4221 786 4233
rect 754 4181 766 4193
rect 694 4167 706 4179
rect 815 4221 827 4233
rect 894 4201 906 4213
rect 1054 4241 1066 4253
rect 1033 4221 1045 4233
rect 973 4201 985 4213
rect 915 4167 927 4179
rect 953 4167 965 4179
rect 1114 4241 1126 4253
rect 1074 4221 1086 4233
rect 1094 4221 1106 4233
rect 1135 4221 1147 4233
rect 1214 4187 1226 4199
rect 1334 4241 1346 4253
rect 1313 4221 1325 4233
rect 1254 4187 1266 4199
rect 1354 4221 1366 4233
rect 1394 4187 1406 4199
rect 1474 4241 1486 4253
rect 1454 4221 1466 4233
rect 1434 4187 1446 4199
rect 1495 4221 1507 4233
rect 1574 4201 1586 4213
rect 1614 4201 1626 4213
rect 1654 4201 1666 4213
rect 1694 4201 1706 4213
rect 1714 4201 1726 4213
rect 1773 4221 1785 4233
rect 1734 4167 1746 4179
rect 1834 4187 1846 4199
rect 1874 4187 1886 4199
rect 1974 4241 1986 4253
rect 1954 4221 1966 4233
rect 1894 4181 1906 4193
rect 2074 4241 2086 4253
rect 1995 4221 2007 4233
rect 2054 4221 2066 4233
rect 2095 4221 2107 4233
rect 2241 4258 2253 4270
rect 2223 4224 2235 4236
rect 2174 4181 2186 4193
rect 2194 4182 2206 4194
rect 2214 4168 2226 4180
rect 2275 4258 2287 4270
rect 2255 4238 2267 4250
rect 2217 4136 2229 4148
rect 2239 4136 2251 4148
rect 2303 4244 2315 4256
rect 2327 4244 2339 4256
rect 2287 4140 2299 4152
rect 2355 4212 2367 4224
rect 2423 4218 2435 4230
rect 2341 4173 2353 4185
rect 2394 4201 2406 4213
rect 2661 4244 2673 4256
rect 2713 4258 2725 4270
rect 2685 4244 2697 4256
rect 2554 4201 2566 4213
rect 2594 4201 2606 4213
rect 2633 4212 2645 4224
rect 2514 4181 2526 4193
rect 2423 4150 2435 4162
rect 2647 4173 2659 4185
rect 2701 4140 2713 4152
rect 2747 4258 2759 4270
rect 2733 4238 2745 4250
rect 2765 4224 2777 4236
rect 2794 4182 2806 4194
rect 2934 4201 2946 4213
rect 2974 4201 2986 4213
rect 2994 4201 3006 4213
rect 2774 4168 2786 4180
rect 2749 4136 2761 4148
rect 2771 4136 2783 4148
rect 2814 4181 2826 4193
rect 2854 4181 2866 4193
rect 3053 4221 3065 4233
rect 3014 4167 3026 4179
rect 3094 4187 3106 4199
rect 3134 4187 3146 4199
rect 3194 4187 3206 4199
rect 3234 4187 3246 4199
rect 3274 4187 3286 4199
rect 3334 4201 3346 4213
rect 3374 4201 3386 4213
rect 3314 4187 3326 4199
rect 3501 4258 3513 4270
rect 3483 4224 3495 4236
rect 3434 4181 3446 4193
rect 3454 4182 3466 4194
rect 3474 4168 3486 4180
rect 3535 4258 3547 4270
rect 3515 4238 3527 4250
rect 3477 4136 3489 4148
rect 3499 4136 3511 4148
rect 3563 4244 3575 4256
rect 3587 4244 3599 4256
rect 3547 4140 3559 4152
rect 3615 4212 3627 4224
rect 3601 4173 3613 4185
rect 3674 4187 3686 4199
rect 3861 4244 3873 4256
rect 3913 4258 3925 4270
rect 3885 4244 3897 4256
rect 3734 4201 3746 4213
rect 3774 4201 3786 4213
rect 3833 4212 3845 4224
rect 3714 4187 3726 4199
rect 3847 4173 3859 4185
rect 3901 4140 3913 4152
rect 3947 4258 3959 4270
rect 3933 4238 3945 4250
rect 3965 4224 3977 4236
rect 3994 4182 4006 4194
rect 4054 4201 4066 4213
rect 4094 4201 4106 4213
rect 3974 4168 3986 4180
rect 3949 4136 3961 4148
rect 3971 4136 3983 4148
rect 4014 4181 4026 4193
rect 4194 4181 4206 4193
rect 4174 4167 4186 4179
rect 4541 4244 4553 4256
rect 4593 4258 4605 4270
rect 4565 4244 4577 4256
rect 4263 4218 4275 4230
rect 4234 4201 4246 4213
rect 4334 4201 4346 4213
rect 4374 4201 4386 4213
rect 4214 4167 4226 4179
rect 4263 4150 4275 4162
rect 4454 4181 4466 4193
rect 4434 4167 4446 4179
rect 4513 4212 4525 4224
rect 4474 4167 4486 4179
rect 4527 4173 4539 4185
rect 4581 4140 4593 4152
rect 4627 4258 4639 4270
rect 4613 4238 4625 4250
rect 4645 4224 4657 4236
rect 4674 4182 4686 4194
rect 4654 4168 4666 4180
rect 4629 4136 4641 4148
rect 4651 4136 4663 4148
rect 4694 4181 4706 4193
rect 34 3981 46 3993
rect 74 3981 86 3993
rect 94 3981 106 3993
rect 134 3981 146 3993
rect 194 3981 206 3993
rect 234 3981 246 3993
rect 314 4001 326 4013
rect 275 3947 287 3959
rect 354 4001 366 4013
rect 334 3967 346 3979
rect 394 4001 406 4013
rect 374 3987 386 3999
rect 534 3981 546 3993
rect 474 3967 486 3979
rect 514 3967 526 3979
rect 574 3981 586 3993
rect 634 4001 646 4013
rect 614 3967 626 3979
rect 673 3947 685 3959
rect 753 3947 765 3959
rect 794 3947 806 3959
rect 814 3947 826 3959
rect 774 3927 786 3939
rect 974 4001 986 4013
rect 855 3947 867 3959
rect 935 3947 947 3959
rect 834 3927 846 3939
rect 1034 4001 1046 4013
rect 994 3967 1006 3979
rect 1014 3967 1026 3979
rect 1154 3987 1166 3999
rect 1073 3947 1085 3959
rect 1213 3947 1225 3959
rect 1274 3987 1286 3999
rect 1254 3947 1266 3959
rect 1234 3927 1246 3939
rect 1334 3947 1346 3959
rect 1375 3947 1387 3959
rect 1434 3947 1446 3959
rect 1354 3927 1366 3939
rect 1534 3981 1546 3993
rect 1475 3947 1487 3959
rect 1454 3927 1466 3939
rect 1574 3981 1586 3993
rect 1733 4018 1745 4030
rect 1634 3967 1646 3979
rect 1674 3967 1686 3979
rect 1734 3981 1746 3993
rect 1774 3967 1786 3979
rect 1854 4001 1866 4013
rect 1815 3947 1827 3959
rect 2014 3987 2026 3999
rect 1874 3967 1886 3979
rect 1894 3967 1906 3979
rect 1934 3967 1946 3979
rect 2054 4001 2066 4013
rect 2034 3967 2046 3979
rect 2134 3987 2146 3999
rect 2093 3947 2105 3959
rect 2194 3981 2206 3993
rect 2234 3981 2246 3993
rect 2274 3947 2286 3959
rect 2403 4018 2415 4030
rect 2374 3967 2386 3979
rect 2315 3947 2327 3959
rect 2294 3927 2306 3939
rect 2474 4001 2486 4013
rect 2510 4004 2522 4016
rect 2550 4004 2562 4016
rect 2590 4004 2602 4016
rect 2403 3950 2415 3962
rect 2674 3987 2686 3999
rect 2717 4032 2729 4044
rect 2739 4032 2751 4044
rect 2714 4000 2726 4012
rect 2694 3986 2706 3998
rect 2723 3944 2735 3956
rect 2755 3930 2767 3942
rect 2741 3910 2753 3922
rect 2787 4028 2799 4040
rect 2841 3995 2853 4007
rect 2894 3987 2906 3999
rect 2855 3956 2867 3968
rect 2803 3924 2815 3936
rect 2775 3910 2787 3922
rect 2827 3924 2839 3936
rect 2974 4001 2986 4013
rect 2954 3967 2966 3979
rect 3134 3981 3146 3993
rect 3054 3967 3066 3979
rect 3013 3947 3025 3959
rect 3094 3967 3106 3979
rect 3254 4001 3266 4013
rect 3174 3981 3186 3993
rect 3294 4001 3306 4013
rect 3274 3987 3286 3999
rect 3355 4018 3367 4030
rect 3354 3981 3366 3993
rect 3314 3967 3326 3979
rect 3534 3987 3546 3999
rect 3434 3967 3446 3979
rect 3474 3967 3486 3979
rect 3587 3995 3599 4007
rect 3573 3956 3585 3968
rect 3641 4028 3653 4040
rect 3601 3924 3613 3936
rect 3625 3924 3637 3936
rect 3689 4032 3701 4044
rect 3711 4032 3723 4044
rect 3673 3930 3685 3942
rect 3653 3910 3665 3922
rect 3714 4000 3726 4012
rect 3834 4001 3846 4013
rect 3734 3986 3746 3998
rect 3754 3987 3766 3999
rect 3705 3944 3717 3956
rect 3687 3910 3699 3922
rect 3874 4001 3886 4013
rect 3854 3987 3866 3999
rect 4095 4018 4107 4030
rect 4094 3981 4106 3993
rect 3894 3967 3906 3979
rect 3934 3967 3946 3979
rect 3994 3967 4006 3979
rect 4034 3967 4046 3979
rect 4054 3967 4066 3979
rect 4174 4001 4186 4013
rect 4154 3967 4166 3979
rect 4314 4001 4326 4013
rect 4213 3947 4225 3959
rect 4275 3947 4287 3959
rect 4394 3987 4406 3999
rect 4334 3967 4346 3979
rect 4447 3995 4459 4007
rect 4433 3956 4445 3968
rect 4501 4028 4513 4040
rect 4461 3924 4473 3936
rect 4485 3924 4497 3936
rect 4549 4032 4561 4044
rect 4571 4032 4583 4044
rect 4533 3930 4545 3942
rect 4513 3910 4525 3922
rect 4574 4000 4586 4012
rect 4594 3986 4606 3998
rect 4614 3987 4626 3999
rect 4654 3987 4666 3999
rect 4565 3944 4577 3956
rect 4547 3910 4559 3922
rect 34 3721 46 3733
rect 74 3721 86 3733
rect 94 3721 106 3733
rect 153 3741 165 3753
rect 114 3687 126 3699
rect 234 3701 246 3713
rect 314 3701 326 3713
rect 294 3687 306 3699
rect 334 3687 346 3699
rect 434 3721 446 3733
rect 394 3707 406 3719
rect 393 3670 405 3682
rect 474 3707 486 3719
rect 514 3707 526 3719
rect 554 3707 566 3719
rect 594 3707 606 3719
rect 674 3721 686 3733
rect 614 3701 626 3713
rect 733 3741 745 3753
rect 694 3687 706 3699
rect 774 3707 786 3719
rect 914 3761 926 3773
rect 893 3741 905 3753
rect 814 3707 826 3719
rect 934 3741 946 3753
rect 974 3701 986 3713
rect 954 3687 966 3699
rect 1074 3761 1086 3773
rect 1054 3741 1066 3753
rect 994 3687 1006 3699
rect 1095 3741 1107 3753
rect 1174 3701 1186 3713
rect 1154 3687 1166 3699
rect 1374 3761 1386 3773
rect 1353 3741 1365 3753
rect 1254 3701 1266 3713
rect 1194 3687 1206 3699
rect 1394 3741 1406 3753
rect 1495 3741 1507 3753
rect 1454 3701 1466 3713
rect 1554 3721 1566 3733
rect 1534 3687 1546 3699
rect 1614 3701 1626 3713
rect 1654 3701 1666 3713
rect 1634 3687 1646 3699
rect 1734 3721 1746 3733
rect 1774 3721 1786 3733
rect 1674 3687 1686 3699
rect 1874 3701 1886 3713
rect 1854 3687 1866 3699
rect 1934 3707 1946 3719
rect 1894 3687 1906 3699
rect 1974 3707 1986 3719
rect 2033 3739 2045 3751
rect 2123 3738 2135 3750
rect 2014 3721 2026 3733
rect 2094 3721 2106 3733
rect 1994 3701 2006 3713
rect 2033 3672 2045 3684
rect 2461 3778 2473 3790
rect 2443 3744 2455 3756
rect 2394 3701 2406 3713
rect 2414 3702 2426 3714
rect 2218 3684 2230 3696
rect 2258 3684 2270 3696
rect 2298 3684 2310 3696
rect 2334 3687 2346 3699
rect 2123 3670 2135 3682
rect 2434 3688 2446 3700
rect 2495 3778 2507 3790
rect 2475 3758 2487 3770
rect 2437 3656 2449 3668
rect 2459 3656 2471 3668
rect 2523 3764 2535 3776
rect 2547 3764 2559 3776
rect 2507 3660 2519 3672
rect 2575 3732 2587 3744
rect 2635 3741 2647 3753
rect 2561 3693 2573 3705
rect 2694 3721 2706 3733
rect 2674 3687 2686 3699
rect 2794 3721 2806 3733
rect 2834 3721 2846 3733
rect 2874 3721 2886 3733
rect 2914 3721 2926 3733
rect 2954 3721 2966 3733
rect 2994 3721 3006 3733
rect 2754 3701 2766 3713
rect 3014 3701 3026 3713
rect 3134 3721 3146 3733
rect 3114 3701 3126 3713
rect 3193 3741 3205 3753
rect 3154 3687 3166 3699
rect 3294 3701 3306 3713
rect 3274 3687 3286 3699
rect 3354 3701 3366 3713
rect 3314 3687 3326 3699
rect 3334 3687 3346 3699
rect 3494 3721 3506 3733
rect 3434 3701 3446 3713
rect 3374 3687 3386 3699
rect 3534 3707 3546 3719
rect 3594 3721 3606 3733
rect 3535 3670 3547 3682
rect 3653 3741 3665 3753
rect 3614 3687 3626 3699
rect 3694 3721 3706 3733
rect 3753 3741 3765 3753
rect 3714 3687 3726 3699
rect 3881 3778 3893 3790
rect 3863 3744 3875 3756
rect 3814 3701 3826 3713
rect 3834 3702 3846 3714
rect 3854 3688 3866 3700
rect 3915 3778 3927 3790
rect 3895 3758 3907 3770
rect 3857 3656 3869 3668
rect 3879 3656 3891 3668
rect 3943 3764 3955 3776
rect 3967 3764 3979 3776
rect 3927 3660 3939 3672
rect 3995 3732 4007 3744
rect 4341 3764 4353 3776
rect 4393 3778 4405 3790
rect 4365 3764 4377 3776
rect 4063 3738 4075 3750
rect 3981 3693 3993 3705
rect 4034 3721 4046 3733
rect 4134 3721 4146 3733
rect 4174 3721 4186 3733
rect 4063 3670 4075 3682
rect 4214 3701 4226 3713
rect 4194 3687 4206 3699
rect 4234 3687 4246 3699
rect 4313 3732 4325 3744
rect 4327 3693 4339 3705
rect 4381 3660 4393 3672
rect 4427 3778 4439 3790
rect 4413 3758 4425 3770
rect 4445 3744 4457 3756
rect 4474 3702 4486 3714
rect 4563 3738 4575 3750
rect 4534 3721 4546 3733
rect 4454 3688 4466 3700
rect 4429 3656 4441 3668
rect 4451 3656 4463 3668
rect 4494 3701 4506 3713
rect 4654 3701 4666 3713
rect 4674 3701 4686 3713
rect 4563 3670 4575 3682
rect 34 3501 46 3513
rect 74 3501 86 3513
rect 114 3507 126 3519
rect 157 3552 169 3564
rect 179 3552 191 3564
rect 154 3520 166 3532
rect 134 3506 146 3518
rect 163 3464 175 3476
rect 195 3450 207 3462
rect 181 3430 193 3442
rect 227 3548 239 3560
rect 281 3515 293 3527
rect 295 3476 307 3488
rect 374 3507 386 3519
rect 243 3444 255 3456
rect 215 3430 227 3442
rect 267 3444 279 3456
rect 414 3501 426 3513
rect 454 3501 466 3513
rect 534 3521 546 3533
rect 495 3467 507 3479
rect 554 3487 566 3499
rect 634 3521 646 3533
rect 595 3467 607 3479
rect 674 3501 686 3513
rect 654 3487 666 3499
rect 714 3501 726 3513
rect 774 3521 786 3533
rect 810 3521 822 3533
rect 754 3487 766 3499
rect 874 3507 886 3519
rect 833 3487 845 3499
rect 973 3467 985 3479
rect 1034 3521 1046 3533
rect 1074 3521 1086 3533
rect 1054 3507 1066 3519
rect 1014 3467 1026 3479
rect 994 3447 1006 3459
rect 1214 3501 1226 3513
rect 1134 3487 1146 3499
rect 1174 3487 1186 3499
rect 1254 3501 1266 3513
rect 1294 3501 1306 3513
rect 1334 3501 1346 3513
rect 1394 3521 1406 3533
rect 1374 3487 1386 3499
rect 1494 3507 1506 3519
rect 1537 3552 1549 3564
rect 1559 3552 1571 3564
rect 1534 3520 1546 3532
rect 1433 3467 1445 3479
rect 1514 3506 1526 3518
rect 1543 3464 1555 3476
rect 1575 3450 1587 3462
rect 1561 3430 1573 3442
rect 1607 3548 1619 3560
rect 1661 3515 1673 3527
rect 1734 3501 1746 3513
rect 1675 3476 1687 3488
rect 1623 3444 1635 3456
rect 1595 3430 1607 3442
rect 1647 3444 1659 3456
rect 1774 3501 1786 3513
rect 1814 3521 1826 3533
rect 1794 3487 1806 3499
rect 1894 3521 1906 3533
rect 1853 3467 1865 3479
rect 2073 3538 2085 3550
rect 1974 3501 1986 3513
rect 2014 3501 2026 3513
rect 2074 3501 2086 3513
rect 2134 3501 2146 3513
rect 2114 3487 2126 3499
rect 2174 3501 2186 3513
rect 2214 3467 2226 3479
rect 2314 3507 2326 3519
rect 2374 3507 2386 3519
rect 2255 3467 2267 3479
rect 2234 3447 2246 3459
rect 2467 3515 2479 3527
rect 2453 3476 2465 3488
rect 2521 3548 2533 3560
rect 2481 3444 2493 3456
rect 2505 3444 2517 3456
rect 2569 3552 2581 3564
rect 2591 3552 2603 3564
rect 2553 3450 2565 3462
rect 2533 3430 2545 3442
rect 2594 3520 2606 3532
rect 2614 3506 2626 3518
rect 2634 3507 2646 3519
rect 2585 3464 2597 3476
rect 2567 3430 2579 3442
rect 2694 3521 2706 3533
rect 2674 3487 2686 3499
rect 2803 3538 2815 3550
rect 2854 3501 2866 3513
rect 2774 3487 2786 3499
rect 2733 3467 2745 3479
rect 2803 3470 2815 3482
rect 2894 3501 2906 3513
rect 2967 3515 2979 3527
rect 2953 3476 2965 3488
rect 3021 3548 3033 3560
rect 2981 3444 2993 3456
rect 3005 3444 3017 3456
rect 3069 3552 3081 3564
rect 3091 3552 3103 3564
rect 3053 3450 3065 3462
rect 3033 3430 3045 3442
rect 3094 3520 3106 3532
rect 3114 3506 3126 3518
rect 3134 3507 3146 3519
rect 3085 3464 3097 3476
rect 3067 3430 3079 3442
rect 3234 3521 3246 3533
rect 3195 3467 3207 3479
rect 3314 3507 3326 3519
rect 3254 3487 3266 3499
rect 3414 3507 3426 3519
rect 3334 3487 3346 3499
rect 3374 3487 3386 3499
rect 3554 3521 3566 3533
rect 3494 3487 3506 3499
rect 3534 3487 3546 3499
rect 3594 3521 3606 3533
rect 3574 3507 3586 3519
rect 3654 3507 3666 3519
rect 3693 3536 3705 3548
rect 3795 3521 3807 3533
rect 3833 3521 3845 3533
rect 3674 3487 3686 3499
rect 3774 3487 3786 3499
rect 3693 3469 3705 3481
rect 3894 3501 3906 3513
rect 3853 3487 3865 3499
rect 3934 3501 3946 3513
rect 3987 3515 3999 3527
rect 3973 3476 3985 3488
rect 4041 3548 4053 3560
rect 4001 3444 4013 3456
rect 4025 3444 4037 3456
rect 4089 3552 4101 3564
rect 4111 3552 4123 3564
rect 4073 3450 4085 3462
rect 4053 3430 4065 3442
rect 4114 3520 4126 3532
rect 4134 3506 4146 3518
rect 4154 3507 4166 3519
rect 4105 3464 4117 3476
rect 4087 3430 4099 3442
rect 4227 3515 4239 3527
rect 4213 3476 4225 3488
rect 4281 3548 4293 3560
rect 4241 3444 4253 3456
rect 4265 3444 4277 3456
rect 4329 3552 4341 3564
rect 4351 3552 4363 3564
rect 4313 3450 4325 3462
rect 4293 3430 4305 3442
rect 4354 3520 4366 3532
rect 4478 3524 4490 3536
rect 4518 3524 4530 3536
rect 4558 3524 4570 3536
rect 4374 3506 4386 3518
rect 4394 3507 4406 3519
rect 4345 3464 4357 3476
rect 4327 3430 4339 3442
rect 4594 3521 4606 3533
rect 4654 3521 4666 3533
rect 4634 3487 4646 3499
rect 4693 3467 4705 3479
rect 101 3298 113 3310
rect 83 3264 95 3276
rect 34 3221 46 3233
rect 54 3222 66 3234
rect 74 3208 86 3220
rect 135 3298 147 3310
rect 115 3278 127 3290
rect 77 3176 89 3188
rect 99 3176 111 3188
rect 163 3284 175 3296
rect 187 3284 199 3296
rect 147 3180 159 3192
rect 215 3252 227 3264
rect 201 3213 213 3225
rect 274 3241 286 3253
rect 353 3241 365 3253
rect 295 3207 307 3219
rect 333 3207 345 3219
rect 394 3227 406 3239
rect 501 3284 513 3296
rect 553 3298 565 3310
rect 525 3284 537 3296
rect 473 3252 485 3264
rect 434 3227 446 3239
rect 487 3213 499 3225
rect 541 3180 553 3192
rect 587 3298 599 3310
rect 573 3278 585 3290
rect 605 3264 617 3276
rect 634 3222 646 3234
rect 715 3261 727 3273
rect 614 3208 626 3220
rect 589 3176 601 3188
rect 611 3176 623 3188
rect 654 3221 666 3233
rect 774 3241 786 3253
rect 814 3241 826 3253
rect 754 3207 766 3219
rect 893 3241 905 3253
rect 835 3207 847 3219
rect 873 3207 885 3219
rect 914 3227 926 3239
rect 1054 3281 1066 3293
rect 1033 3261 1045 3273
rect 954 3227 966 3239
rect 1074 3261 1086 3273
rect 1214 3281 1226 3293
rect 1194 3261 1206 3273
rect 1174 3241 1186 3253
rect 1134 3227 1146 3239
rect 1133 3190 1145 3202
rect 1235 3261 1247 3273
rect 1294 3241 1306 3253
rect 1353 3261 1365 3273
rect 1314 3207 1326 3219
rect 1394 3227 1406 3239
rect 1515 3259 1527 3271
rect 1534 3241 1546 3253
rect 1434 3227 1446 3239
rect 1515 3192 1527 3204
rect 1554 3221 1566 3233
rect 1594 3227 1606 3239
rect 1654 3241 1666 3253
rect 1634 3227 1646 3239
rect 1713 3261 1725 3273
rect 1775 3261 1787 3273
rect 1674 3207 1686 3219
rect 1834 3241 1846 3253
rect 1814 3207 1826 3219
rect 1854 3227 1866 3239
rect 1934 3241 1946 3253
rect 1894 3227 1906 3239
rect 1993 3261 2005 3273
rect 2055 3261 2067 3273
rect 1954 3207 1966 3219
rect 2114 3241 2126 3253
rect 2094 3207 2106 3219
rect 2194 3241 2206 3253
rect 2134 3221 2146 3233
rect 2253 3261 2265 3273
rect 2214 3207 2226 3219
rect 2334 3221 2346 3233
rect 2354 3227 2366 3239
rect 2481 3284 2493 3296
rect 2533 3298 2545 3310
rect 2505 3284 2517 3296
rect 2453 3252 2465 3264
rect 2394 3227 2406 3239
rect 2467 3213 2479 3225
rect 2521 3180 2533 3192
rect 2567 3298 2579 3310
rect 2553 3278 2565 3290
rect 2585 3264 2597 3276
rect 2614 3222 2626 3234
rect 2801 3284 2813 3296
rect 2853 3298 2865 3310
rect 2825 3284 2837 3296
rect 2703 3258 2715 3270
rect 2674 3241 2686 3253
rect 2594 3208 2606 3220
rect 2569 3176 2581 3188
rect 2591 3176 2603 3188
rect 2634 3221 2646 3233
rect 2773 3252 2785 3264
rect 2703 3190 2715 3202
rect 2787 3213 2799 3225
rect 2841 3180 2853 3192
rect 2887 3298 2899 3310
rect 2873 3278 2885 3290
rect 2905 3264 2917 3276
rect 2934 3222 2946 3234
rect 3015 3261 3027 3273
rect 2914 3208 2926 3220
rect 2889 3176 2901 3188
rect 2911 3176 2923 3188
rect 2954 3221 2966 3233
rect 3115 3261 3127 3273
rect 3074 3241 3086 3253
rect 3054 3207 3066 3219
rect 3174 3241 3186 3253
rect 3194 3241 3206 3253
rect 3154 3207 3166 3219
rect 3253 3261 3265 3273
rect 3315 3261 3327 3273
rect 3214 3207 3226 3219
rect 3374 3241 3386 3253
rect 3394 3241 3406 3253
rect 3354 3207 3366 3219
rect 3453 3261 3465 3273
rect 3414 3207 3426 3219
rect 3494 3227 3506 3239
rect 3534 3227 3546 3239
rect 3574 3227 3586 3239
rect 3614 3227 3626 3239
rect 3654 3227 3666 3239
rect 3694 3227 3706 3239
rect 3734 3227 3746 3239
rect 3843 3258 3855 3270
rect 3814 3241 3826 3253
rect 3774 3227 3786 3239
rect 3914 3227 3926 3239
rect 3994 3241 4006 3253
rect 4083 3258 4095 3270
rect 4034 3241 4046 3253
rect 4054 3241 4066 3253
rect 3954 3227 3966 3239
rect 3843 3190 3855 3202
rect 4215 3261 4227 3273
rect 4174 3221 4186 3233
rect 4083 3190 4095 3202
rect 4274 3241 4286 3253
rect 4254 3207 4266 3219
rect 4354 3241 4366 3253
rect 4334 3221 4346 3233
rect 4413 3261 4425 3273
rect 4374 3207 4386 3219
rect 4474 3227 4486 3239
rect 4514 3227 4526 3239
rect 4621 3298 4633 3310
rect 4603 3264 4615 3276
rect 4554 3221 4566 3233
rect 4574 3222 4586 3234
rect 4594 3208 4606 3220
rect 4655 3298 4667 3310
rect 4635 3278 4647 3290
rect 4597 3176 4609 3188
rect 4619 3176 4631 3188
rect 4683 3284 4695 3296
rect 4707 3284 4719 3296
rect 4667 3180 4679 3192
rect 4735 3252 4747 3264
rect 4721 3213 4733 3225
rect 55 3041 67 3053
rect 93 3041 105 3053
rect 34 3007 46 3019
rect 173 3058 185 3070
rect 113 3007 125 3019
rect 174 3021 186 3033
rect 214 3007 226 3019
rect 267 3035 279 3047
rect 253 2996 265 3008
rect 321 3068 333 3080
rect 281 2964 293 2976
rect 305 2964 317 2976
rect 369 3072 381 3084
rect 391 3072 403 3084
rect 353 2970 365 2982
rect 333 2950 345 2962
rect 394 3040 406 3052
rect 414 3026 426 3038
rect 434 3027 446 3039
rect 385 2984 397 2996
rect 367 2950 379 2962
rect 494 3041 506 3053
rect 474 3007 486 3019
rect 574 3021 586 3033
rect 533 2987 545 2999
rect 614 3021 626 3033
rect 674 3021 686 3033
rect 714 3021 726 3033
rect 814 3021 826 3033
rect 754 3007 766 3019
rect 794 3007 806 3019
rect 854 3021 866 3033
rect 954 3041 966 3053
rect 915 2987 927 2999
rect 974 3007 986 3019
rect 1054 3041 1066 3053
rect 1015 2987 1027 2999
rect 1074 3007 1086 3019
rect 1114 3007 1126 3019
rect 1154 3007 1166 3019
rect 1234 3041 1246 3053
rect 1195 2987 1207 2999
rect 1274 3021 1286 3033
rect 1254 3007 1266 3019
rect 1394 3041 1406 3053
rect 1314 3021 1326 3033
rect 1414 3021 1426 3033
rect 1454 3021 1466 3033
rect 1494 3021 1506 3033
rect 1534 3021 1546 3033
rect 1603 3058 1615 3070
rect 1674 3041 1686 3053
rect 1574 3007 1586 3019
rect 1654 3007 1666 3019
rect 1603 2990 1615 3002
rect 1774 3041 1786 3053
rect 1754 3007 1766 3019
rect 1713 2987 1725 2999
rect 1934 3041 1946 3053
rect 1854 3007 1866 3019
rect 1813 2987 1825 2999
rect 1894 3007 1906 3019
rect 1974 3041 1986 3053
rect 1954 3027 1966 3039
rect 2034 3027 2046 3039
rect 2114 3041 2126 3053
rect 2094 3007 2106 3019
rect 2294 3021 2306 3033
rect 2194 3007 2206 3019
rect 2153 2987 2165 2999
rect 2234 3007 2246 3019
rect 2334 3021 2346 3033
rect 2374 3041 2386 3053
rect 2354 3007 2366 3019
rect 2454 3027 2466 3039
rect 2413 2987 2425 2999
rect 2534 3041 2546 3053
rect 2514 3007 2526 3019
rect 2643 3058 2655 3070
rect 2694 3021 2706 3033
rect 2614 3007 2626 3019
rect 2573 2987 2585 2999
rect 2643 2990 2655 3002
rect 2734 3021 2746 3033
rect 2794 3027 2806 3039
rect 2837 3072 2849 3084
rect 2859 3072 2871 3084
rect 2834 3040 2846 3052
rect 2814 3026 2826 3038
rect 2843 2984 2855 2996
rect 2875 2970 2887 2982
rect 2861 2950 2873 2962
rect 2907 3068 2919 3080
rect 2961 3035 2973 3047
rect 3134 3041 3146 3053
rect 2975 2996 2987 3008
rect 3034 3007 3046 3019
rect 3074 3007 3086 3019
rect 3174 3041 3186 3053
rect 3154 3027 3166 3039
rect 3294 3027 3306 3039
rect 3337 3072 3349 3084
rect 3359 3072 3371 3084
rect 3334 3040 3346 3052
rect 3194 3007 3206 3019
rect 3234 3007 3246 3019
rect 3314 3026 3326 3038
rect 2923 2964 2935 2976
rect 2895 2950 2907 2962
rect 2947 2964 2959 2976
rect 3343 2984 3355 2996
rect 3375 2970 3387 2982
rect 3361 2950 3373 2962
rect 3407 3068 3419 3080
rect 3461 3035 3473 3047
rect 3534 3027 3546 3039
rect 3577 3072 3589 3084
rect 3599 3072 3611 3084
rect 3574 3040 3586 3052
rect 3475 2996 3487 3008
rect 3554 3026 3566 3038
rect 3423 2964 3435 2976
rect 3395 2950 3407 2962
rect 3447 2964 3459 2976
rect 3583 2984 3595 2996
rect 3615 2970 3627 2982
rect 3601 2950 3613 2962
rect 3647 3068 3659 3080
rect 3701 3035 3713 3047
rect 3715 2996 3727 3008
rect 3754 3007 3766 3019
rect 3794 3007 3806 3019
rect 3894 3041 3906 3053
rect 3855 2987 3867 2999
rect 3663 2964 3675 2976
rect 3635 2950 3647 2962
rect 3687 2964 3699 2976
rect 3914 3007 3926 3019
rect 3994 3041 4006 3053
rect 3955 2987 3967 2999
rect 4054 3041 4066 3053
rect 4014 3007 4026 3019
rect 4034 3007 4046 3019
rect 4154 3041 4166 3053
rect 4134 3007 4146 3019
rect 4093 2987 4105 2999
rect 4234 3027 4246 3039
rect 4193 2987 4205 2999
rect 4294 2987 4306 2999
rect 4427 3035 4439 3047
rect 4335 2987 4347 2999
rect 4314 2967 4326 2979
rect 4413 2996 4425 3008
rect 4481 3068 4493 3080
rect 4441 2964 4453 2976
rect 4465 2964 4477 2976
rect 4529 3072 4541 3084
rect 4551 3072 4563 3084
rect 4513 2970 4525 2982
rect 4493 2950 4505 2962
rect 4554 3040 4566 3052
rect 4574 3026 4586 3038
rect 4594 3027 4606 3039
rect 4545 2984 4557 2996
rect 4527 2950 4539 2962
rect 4654 3041 4666 3053
rect 4634 3007 4646 3019
rect 4693 2987 4705 2999
rect 95 2781 107 2793
rect 54 2741 66 2753
rect 154 2761 166 2773
rect 175 2761 187 2773
rect 134 2727 146 2739
rect 254 2761 266 2773
rect 195 2727 207 2739
rect 233 2727 245 2739
rect 294 2747 306 2759
rect 374 2761 386 2773
rect 334 2747 346 2759
rect 414 2747 426 2759
rect 495 2781 507 2793
rect 415 2710 427 2722
rect 554 2761 566 2773
rect 534 2727 546 2739
rect 574 2747 586 2759
rect 614 2747 626 2759
rect 774 2747 786 2759
rect 694 2727 706 2739
rect 754 2727 766 2739
rect 854 2761 866 2773
rect 814 2747 826 2759
rect 894 2747 906 2759
rect 975 2781 987 2793
rect 895 2710 907 2722
rect 1034 2761 1046 2773
rect 1014 2727 1026 2739
rect 1054 2747 1066 2759
rect 1281 2804 1293 2816
rect 1333 2818 1345 2830
rect 1305 2804 1317 2816
rect 1155 2781 1167 2793
rect 1094 2747 1106 2759
rect 1214 2761 1226 2773
rect 1253 2772 1265 2784
rect 1194 2727 1206 2739
rect 1267 2733 1279 2745
rect 1321 2700 1333 2712
rect 1367 2818 1379 2830
rect 1353 2798 1365 2810
rect 1385 2784 1397 2796
rect 1414 2742 1426 2754
rect 1505 2778 1517 2790
rect 1534 2761 1546 2773
rect 1394 2728 1406 2740
rect 1369 2696 1381 2708
rect 1391 2696 1403 2708
rect 1434 2741 1446 2753
rect 1505 2710 1517 2722
rect 1641 2818 1653 2830
rect 1623 2784 1635 2796
rect 1574 2741 1586 2753
rect 1594 2742 1606 2754
rect 1614 2728 1626 2740
rect 1675 2818 1687 2830
rect 1655 2798 1667 2810
rect 1617 2696 1629 2708
rect 1639 2696 1651 2708
rect 1703 2804 1715 2816
rect 1727 2804 1739 2816
rect 1687 2700 1699 2712
rect 1755 2772 1767 2784
rect 1741 2733 1753 2745
rect 1794 2761 1806 2773
rect 1853 2781 1865 2793
rect 1814 2727 1826 2739
rect 1954 2761 1966 2773
rect 1894 2741 1906 2753
rect 2033 2761 2045 2773
rect 2094 2761 2106 2773
rect 2134 2761 2146 2773
rect 2174 2761 2186 2773
rect 2214 2761 2226 2773
rect 2254 2761 2266 2773
rect 2294 2761 2306 2773
rect 1974 2727 1986 2739
rect 2010 2727 2022 2739
rect 2394 2761 2406 2773
rect 2434 2761 2446 2773
rect 2314 2741 2326 2753
rect 2514 2761 2526 2773
rect 2454 2741 2466 2753
rect 2554 2747 2566 2759
rect 2614 2761 2626 2773
rect 2555 2710 2567 2722
rect 2673 2781 2685 2793
rect 2634 2727 2646 2739
rect 2714 2761 2726 2773
rect 2773 2781 2785 2793
rect 2734 2727 2746 2739
rect 2814 2747 2826 2759
rect 2854 2747 2866 2759
rect 2981 2818 2993 2830
rect 2963 2784 2975 2796
rect 2914 2741 2926 2753
rect 2934 2742 2946 2754
rect 2954 2728 2966 2740
rect 3015 2818 3027 2830
rect 2995 2798 3007 2810
rect 2957 2696 2969 2708
rect 2979 2696 2991 2708
rect 3043 2804 3055 2816
rect 3067 2804 3079 2816
rect 3027 2700 3039 2712
rect 3095 2772 3107 2784
rect 3081 2733 3093 2745
rect 3221 2818 3233 2830
rect 3203 2784 3215 2796
rect 3154 2741 3166 2753
rect 3174 2742 3186 2754
rect 3194 2728 3206 2740
rect 3255 2818 3267 2830
rect 3235 2798 3247 2810
rect 3197 2696 3209 2708
rect 3219 2696 3231 2708
rect 3283 2804 3295 2816
rect 3307 2804 3319 2816
rect 3267 2700 3279 2712
rect 3335 2772 3347 2784
rect 3321 2733 3333 2745
rect 3454 2761 3466 2773
rect 3494 2761 3506 2773
rect 3414 2741 3426 2753
rect 3661 2818 3673 2830
rect 3643 2784 3655 2796
rect 3594 2741 3606 2753
rect 3614 2742 3626 2754
rect 3554 2727 3566 2739
rect 3634 2728 3646 2740
rect 3695 2818 3707 2830
rect 3675 2798 3687 2810
rect 3637 2696 3649 2708
rect 3659 2696 3671 2708
rect 3723 2804 3735 2816
rect 3747 2804 3759 2816
rect 3707 2700 3719 2712
rect 3775 2772 3787 2784
rect 3761 2733 3773 2745
rect 3834 2761 3846 2773
rect 3913 2761 3925 2773
rect 3954 2761 3966 2773
rect 3994 2761 4006 2773
rect 4014 2761 4026 2773
rect 3855 2727 3867 2739
rect 3893 2727 3905 2739
rect 4073 2781 4085 2793
rect 4135 2781 4147 2793
rect 4034 2727 4046 2739
rect 4194 2761 4206 2773
rect 4214 2761 4226 2773
rect 4254 2761 4266 2773
rect 4174 2727 4186 2739
rect 4381 2818 4393 2830
rect 4363 2784 4375 2796
rect 4314 2741 4326 2753
rect 4334 2742 4346 2754
rect 4354 2728 4366 2740
rect 4415 2818 4427 2830
rect 4395 2798 4407 2810
rect 4357 2696 4369 2708
rect 4379 2696 4391 2708
rect 4443 2804 4455 2816
rect 4467 2804 4479 2816
rect 4427 2700 4439 2712
rect 4495 2772 4507 2784
rect 4481 2733 4493 2745
rect 4534 2761 4546 2773
rect 4593 2781 4605 2793
rect 4554 2727 4566 2739
rect 4634 2747 4646 2759
rect 4674 2747 4686 2759
rect 14 2507 26 2519
rect 114 2561 126 2573
rect 154 2561 166 2573
rect 134 2547 146 2559
rect 55 2507 67 2519
rect 34 2487 46 2499
rect 313 2578 325 2590
rect 254 2547 266 2559
rect 314 2541 326 2553
rect 414 2561 426 2573
rect 354 2527 366 2539
rect 454 2561 466 2573
rect 434 2547 446 2559
rect 513 2507 525 2519
rect 634 2561 646 2573
rect 554 2507 566 2519
rect 595 2507 607 2519
rect 534 2487 546 2499
rect 714 2561 726 2573
rect 654 2527 666 2539
rect 754 2541 766 2553
rect 794 2541 806 2553
rect 853 2507 865 2519
rect 974 2561 986 2573
rect 894 2507 906 2519
rect 935 2507 947 2519
rect 874 2487 886 2499
rect 1014 2541 1026 2553
rect 994 2527 1006 2539
rect 1054 2541 1066 2553
rect 1133 2507 1145 2519
rect 1234 2547 1246 2559
rect 1174 2507 1186 2519
rect 1154 2487 1166 2499
rect 1314 2561 1326 2573
rect 1275 2507 1287 2519
rect 1354 2541 1366 2553
rect 1334 2527 1346 2539
rect 1434 2561 1446 2573
rect 1394 2541 1406 2553
rect 1514 2541 1526 2553
rect 1554 2541 1566 2553
rect 1594 2547 1606 2559
rect 1637 2592 1649 2604
rect 1659 2592 1671 2604
rect 1634 2560 1646 2572
rect 1614 2546 1626 2558
rect 1643 2504 1655 2516
rect 1675 2490 1687 2502
rect 1661 2470 1673 2482
rect 1707 2588 1719 2600
rect 1761 2555 1773 2567
rect 1814 2541 1826 2553
rect 1775 2516 1787 2528
rect 1723 2484 1735 2496
rect 1695 2470 1707 2482
rect 1747 2484 1759 2496
rect 1854 2541 1866 2553
rect 1894 2541 1906 2553
rect 1934 2541 1946 2553
rect 1974 2507 1986 2519
rect 2194 2547 2206 2559
rect 2074 2527 2086 2539
rect 2015 2507 2027 2519
rect 1994 2487 2006 2499
rect 2114 2527 2126 2539
rect 2334 2547 2346 2559
rect 2234 2527 2246 2539
rect 2274 2527 2286 2539
rect 2414 2561 2426 2573
rect 2375 2507 2387 2519
rect 2575 2578 2587 2590
rect 2574 2541 2586 2553
rect 2434 2527 2446 2539
rect 2454 2527 2466 2539
rect 2494 2527 2506 2539
rect 2534 2527 2546 2539
rect 2654 2561 2666 2573
rect 2634 2527 2646 2539
rect 2754 2541 2766 2553
rect 2693 2507 2705 2519
rect 2794 2541 2806 2553
rect 2814 2547 2826 2559
rect 2853 2576 2865 2588
rect 2914 2541 2926 2553
rect 2834 2527 2846 2539
rect 2853 2509 2865 2521
rect 2954 2541 2966 2553
rect 3023 2578 3035 2590
rect 3094 2561 3106 2573
rect 2994 2527 3006 2539
rect 3074 2527 3086 2539
rect 3023 2510 3035 2522
rect 3205 2578 3217 2590
rect 3274 2541 3286 2553
rect 3234 2527 3246 2539
rect 3133 2507 3145 2519
rect 3205 2510 3217 2522
rect 3314 2541 3326 2553
rect 3355 2561 3367 2573
rect 3393 2561 3405 2573
rect 3335 2527 3347 2539
rect 3483 2578 3495 2590
rect 3565 2578 3577 2590
rect 3414 2527 3426 2539
rect 3454 2527 3466 2539
rect 3634 2547 3646 2559
rect 3677 2592 3689 2604
rect 3699 2592 3711 2604
rect 3674 2560 3686 2572
rect 3594 2527 3606 2539
rect 3483 2510 3495 2522
rect 3565 2510 3577 2522
rect 3654 2546 3666 2558
rect 3683 2504 3695 2516
rect 3715 2490 3727 2502
rect 3701 2470 3713 2482
rect 3747 2588 3759 2600
rect 3801 2555 3813 2567
rect 3815 2516 3827 2528
rect 3894 2561 3906 2573
rect 3934 2561 3946 2573
rect 3914 2547 3926 2559
rect 4054 2561 4066 2573
rect 4090 2564 4102 2576
rect 4130 2564 4142 2576
rect 4170 2564 4182 2576
rect 3954 2527 3966 2539
rect 3994 2527 4006 2539
rect 4254 2547 4266 2559
rect 4297 2592 4309 2604
rect 4319 2592 4331 2604
rect 4294 2560 4306 2572
rect 4274 2546 4286 2558
rect 3763 2484 3775 2496
rect 3735 2470 3747 2482
rect 3787 2484 3799 2496
rect 4303 2504 4315 2516
rect 4335 2490 4347 2502
rect 4321 2470 4333 2482
rect 4367 2588 4379 2600
rect 4421 2555 4433 2567
rect 4494 2561 4506 2573
rect 4435 2516 4447 2528
rect 4474 2527 4486 2539
rect 4574 2541 4586 2553
rect 4533 2507 4545 2519
rect 4383 2484 4395 2496
rect 4355 2470 4367 2482
rect 4407 2484 4419 2496
rect 4614 2541 4626 2553
rect 4654 2541 4666 2553
rect 4694 2541 4706 2553
rect 74 2321 86 2333
rect 53 2301 65 2313
rect 94 2301 106 2313
rect 135 2301 147 2313
rect 194 2281 206 2293
rect 214 2281 226 2293
rect 174 2247 186 2259
rect 334 2321 346 2333
rect 273 2301 285 2313
rect 314 2301 326 2313
rect 234 2247 246 2259
rect 355 2301 367 2313
rect 434 2261 446 2273
rect 414 2247 426 2259
rect 514 2281 526 2293
rect 454 2247 466 2259
rect 573 2301 585 2313
rect 534 2247 546 2259
rect 674 2261 686 2273
rect 654 2247 666 2259
rect 714 2261 726 2273
rect 694 2247 706 2259
rect 854 2281 866 2293
rect 814 2267 826 2279
rect 813 2230 825 2242
rect 874 2267 886 2279
rect 954 2281 966 2293
rect 914 2267 926 2279
rect 994 2267 1006 2279
rect 1075 2301 1087 2313
rect 995 2230 1007 2242
rect 1175 2301 1187 2313
rect 1134 2281 1146 2293
rect 1114 2247 1126 2259
rect 1234 2281 1246 2293
rect 1214 2247 1226 2259
rect 1341 2338 1353 2350
rect 1323 2304 1335 2316
rect 1274 2261 1286 2273
rect 1294 2262 1306 2274
rect 1314 2248 1326 2260
rect 1375 2338 1387 2350
rect 1355 2318 1367 2330
rect 1317 2216 1329 2228
rect 1339 2216 1351 2228
rect 1403 2324 1415 2336
rect 1427 2324 1439 2336
rect 1387 2220 1399 2232
rect 1455 2292 1467 2304
rect 1515 2301 1527 2313
rect 1441 2253 1453 2265
rect 1574 2281 1586 2293
rect 1554 2247 1566 2259
rect 1681 2338 1693 2350
rect 1663 2304 1675 2316
rect 1614 2261 1626 2273
rect 1634 2262 1646 2274
rect 1654 2248 1666 2260
rect 1715 2338 1727 2350
rect 1695 2318 1707 2330
rect 1657 2216 1669 2228
rect 1679 2216 1691 2228
rect 1743 2324 1755 2336
rect 1767 2324 1779 2336
rect 1727 2220 1739 2232
rect 1795 2292 1807 2304
rect 1781 2253 1793 2265
rect 1954 2281 1966 2293
rect 1874 2261 1886 2273
rect 1934 2261 1946 2273
rect 2013 2301 2025 2313
rect 1974 2247 1986 2259
rect 2141 2338 2153 2350
rect 2123 2304 2135 2316
rect 2074 2261 2086 2273
rect 2094 2262 2106 2274
rect 2114 2248 2126 2260
rect 2175 2338 2187 2350
rect 2155 2318 2167 2330
rect 2117 2216 2129 2228
rect 2139 2216 2151 2228
rect 2203 2324 2215 2336
rect 2227 2324 2239 2336
rect 2187 2220 2199 2232
rect 2255 2292 2267 2304
rect 2241 2253 2253 2265
rect 2354 2261 2366 2273
rect 2334 2247 2346 2259
rect 2514 2321 2526 2333
rect 2494 2301 2506 2313
rect 2454 2261 2466 2273
rect 2374 2247 2386 2259
rect 2434 2247 2446 2259
rect 2474 2247 2486 2259
rect 2535 2301 2547 2313
rect 2594 2281 2606 2293
rect 2741 2324 2753 2336
rect 2793 2338 2805 2350
rect 2765 2324 2777 2336
rect 2634 2267 2646 2279
rect 2635 2230 2647 2242
rect 2713 2292 2725 2304
rect 2727 2253 2739 2265
rect 2781 2220 2793 2232
rect 2827 2338 2839 2350
rect 2813 2318 2825 2330
rect 2845 2304 2857 2316
rect 2874 2262 2886 2274
rect 2955 2301 2967 2313
rect 2854 2248 2866 2260
rect 2829 2216 2841 2228
rect 2851 2216 2863 2228
rect 2894 2261 2906 2273
rect 3055 2301 3067 2313
rect 3014 2281 3026 2293
rect 2994 2247 3006 2259
rect 3114 2281 3126 2293
rect 3134 2281 3146 2293
rect 3094 2247 3106 2259
rect 3281 2324 3293 2336
rect 3333 2338 3345 2350
rect 3305 2324 3317 2336
rect 3193 2301 3205 2313
rect 3154 2247 3166 2259
rect 3253 2292 3265 2304
rect 3267 2253 3279 2265
rect 3321 2220 3333 2232
rect 3367 2338 3379 2350
rect 3353 2318 3365 2330
rect 3385 2304 3397 2316
rect 3414 2262 3426 2274
rect 3495 2301 3507 2313
rect 3394 2248 3406 2260
rect 3369 2216 3381 2228
rect 3391 2216 3403 2228
rect 3434 2261 3446 2273
rect 3554 2281 3566 2293
rect 3594 2281 3606 2293
rect 3634 2281 3646 2293
rect 3534 2247 3546 2259
rect 3693 2299 3705 2311
rect 3674 2281 3686 2293
rect 3654 2261 3666 2273
rect 3774 2267 3786 2279
rect 3854 2281 3866 2293
rect 3814 2267 3826 2279
rect 3693 2232 3705 2244
rect 3933 2281 3945 2293
rect 3974 2281 3986 2293
rect 3875 2247 3887 2259
rect 3913 2247 3925 2259
rect 4053 2281 4065 2293
rect 3995 2247 4007 2259
rect 4033 2247 4045 2259
rect 4161 2338 4173 2350
rect 4143 2304 4155 2316
rect 4094 2261 4106 2273
rect 4114 2262 4126 2274
rect 4134 2248 4146 2260
rect 4195 2338 4207 2350
rect 4175 2318 4187 2330
rect 4137 2216 4149 2228
rect 4159 2216 4171 2228
rect 4223 2324 4235 2336
rect 4247 2324 4259 2336
rect 4207 2220 4219 2232
rect 4361 2324 4373 2336
rect 4413 2338 4425 2350
rect 4385 2324 4397 2336
rect 4275 2292 4287 2304
rect 4261 2253 4273 2265
rect 4333 2292 4345 2304
rect 4347 2253 4359 2265
rect 4401 2220 4413 2232
rect 4447 2338 4459 2350
rect 4433 2318 4445 2330
rect 4465 2304 4477 2316
rect 4494 2262 4506 2274
rect 4554 2281 4566 2293
rect 4474 2248 4486 2260
rect 4449 2216 4461 2228
rect 4471 2216 4483 2228
rect 4514 2261 4526 2273
rect 4613 2301 4625 2313
rect 4574 2247 4586 2259
rect 4654 2267 4666 2279
rect 4694 2267 4706 2279
rect 45 2098 57 2110
rect 74 2047 86 2059
rect 45 2030 57 2042
rect 154 2081 166 2093
rect 115 2027 127 2039
rect 174 2047 186 2059
rect 233 2027 245 2039
rect 294 2081 306 2093
rect 334 2081 346 2093
rect 394 2081 406 2093
rect 314 2067 326 2079
rect 274 2027 286 2039
rect 254 2007 266 2019
rect 434 2081 446 2093
rect 414 2067 426 2079
rect 494 2027 506 2039
rect 535 2027 547 2039
rect 594 2027 606 2039
rect 514 2007 526 2019
rect 694 2081 706 2093
rect 734 2081 746 2093
rect 714 2067 726 2079
rect 635 2027 647 2039
rect 614 2007 626 2019
rect 854 2081 866 2093
rect 815 2027 827 2039
rect 874 2047 886 2059
rect 894 2027 906 2039
rect 935 2027 947 2039
rect 994 2027 1006 2039
rect 914 2007 926 2019
rect 1035 2027 1047 2039
rect 1094 2027 1106 2039
rect 1014 2007 1026 2019
rect 1194 2081 1206 2093
rect 1234 2081 1246 2093
rect 1214 2067 1226 2079
rect 1135 2027 1147 2039
rect 1114 2007 1126 2019
rect 1394 2061 1406 2073
rect 1294 2047 1306 2059
rect 1334 2047 1346 2059
rect 1434 2061 1446 2073
rect 1474 2061 1486 2073
rect 1514 2061 1526 2073
rect 1534 2061 1546 2073
rect 1574 2061 1586 2073
rect 1674 2081 1686 2093
rect 1635 2027 1647 2039
rect 1714 2081 1726 2093
rect 1694 2047 1706 2059
rect 1754 2081 1766 2093
rect 1734 2067 1746 2079
rect 1814 2047 1826 2059
rect 1854 2047 1866 2059
rect 1954 2081 1966 2093
rect 1915 2027 1927 2039
rect 2014 2081 2026 2093
rect 1974 2047 1986 2059
rect 1994 2047 2006 2059
rect 2154 2081 2166 2093
rect 2053 2027 2065 2039
rect 2115 2027 2127 2039
rect 2238 2084 2250 2096
rect 2278 2084 2290 2096
rect 2318 2084 2330 2096
rect 2174 2047 2186 2059
rect 2354 2081 2366 2093
rect 2513 2098 2525 2110
rect 2394 2061 2406 2073
rect 2434 2061 2446 2073
rect 2514 2061 2526 2073
rect 2574 2067 2586 2079
rect 2554 2047 2566 2059
rect 2613 2096 2625 2108
rect 2694 2061 2706 2073
rect 2594 2047 2606 2059
rect 2613 2029 2625 2041
rect 2734 2061 2746 2073
rect 2754 2061 2766 2073
rect 2794 2061 2806 2073
rect 2854 2067 2866 2079
rect 2897 2112 2909 2124
rect 2919 2112 2931 2124
rect 2894 2080 2906 2092
rect 2874 2066 2886 2078
rect 2903 2024 2915 2036
rect 2935 2010 2947 2022
rect 2921 1990 2933 2002
rect 2967 2108 2979 2120
rect 3021 2075 3033 2087
rect 3035 2036 3047 2048
rect 3114 2081 3126 2093
rect 3154 2081 3166 2093
rect 3134 2067 3146 2079
rect 3295 2081 3307 2093
rect 3333 2081 3345 2093
rect 3174 2047 3186 2059
rect 3214 2047 3226 2059
rect 3274 2047 3286 2059
rect 3394 2067 3406 2079
rect 3437 2112 3449 2124
rect 3459 2112 3471 2124
rect 3434 2080 3446 2092
rect 3353 2047 3365 2059
rect 3414 2066 3426 2078
rect 2983 2004 2995 2016
rect 2955 1990 2967 2002
rect 3007 2004 3019 2016
rect 3443 2024 3455 2036
rect 3475 2010 3487 2022
rect 3461 1990 3473 2002
rect 3507 2108 3519 2120
rect 3561 2075 3573 2087
rect 3634 2081 3646 2093
rect 3575 2036 3587 2048
rect 3614 2047 3626 2059
rect 3734 2067 3746 2079
rect 3777 2112 3789 2124
rect 3799 2112 3811 2124
rect 3774 2080 3786 2092
rect 3673 2027 3685 2039
rect 3523 2004 3535 2016
rect 3495 1990 3507 2002
rect 3547 2004 3559 2016
rect 3754 2066 3766 2078
rect 3783 2024 3795 2036
rect 3815 2010 3827 2022
rect 3801 1990 3813 2002
rect 3847 2108 3859 2120
rect 3901 2075 3913 2087
rect 3915 2036 3927 2048
rect 3987 2075 3999 2087
rect 3973 2036 3985 2048
rect 3863 2004 3875 2016
rect 3835 1990 3847 2002
rect 3887 2004 3899 2016
rect 4041 2108 4053 2120
rect 4001 2004 4013 2016
rect 4025 2004 4037 2016
rect 4089 2112 4101 2124
rect 4111 2112 4123 2124
rect 4073 2010 4085 2022
rect 4053 1990 4065 2002
rect 4114 2080 4126 2092
rect 4134 2066 4146 2078
rect 4154 2067 4166 2079
rect 4105 2024 4117 2036
rect 4087 1990 4099 2002
rect 4235 2081 4247 2093
rect 4273 2081 4285 2093
rect 4214 2047 4226 2059
rect 4314 2067 4326 2079
rect 4293 2047 4305 2059
rect 4394 2047 4406 2059
rect 4434 2047 4446 2059
rect 4474 2047 4486 2059
rect 4514 2047 4526 2059
rect 4567 2075 4579 2087
rect 4553 2036 4565 2048
rect 4621 2108 4633 2120
rect 4581 2004 4593 2016
rect 4605 2004 4617 2016
rect 4669 2112 4681 2124
rect 4691 2112 4703 2124
rect 4653 2010 4665 2022
rect 4633 1990 4645 2002
rect 4694 2080 4706 2092
rect 4714 2066 4726 2078
rect 4734 2067 4746 2079
rect 4685 2024 4697 2036
rect 4667 1990 4679 2002
rect 34 1801 46 1813
rect 113 1801 125 1813
rect 134 1801 146 1813
rect 55 1767 67 1779
rect 93 1767 105 1779
rect 193 1821 205 1833
rect 154 1767 166 1779
rect 234 1787 246 1799
rect 374 1841 386 1853
rect 353 1821 365 1833
rect 274 1787 286 1799
rect 394 1821 406 1833
rect 415 1801 427 1813
rect 494 1801 506 1813
rect 534 1801 546 1813
rect 435 1767 447 1779
rect 473 1767 485 1779
rect 574 1787 586 1799
rect 575 1750 587 1762
rect 723 1818 735 1830
rect 795 1821 807 1833
rect 694 1801 706 1813
rect 674 1767 686 1779
rect 723 1750 735 1762
rect 854 1801 866 1813
rect 874 1801 886 1813
rect 834 1767 846 1779
rect 994 1841 1006 1853
rect 933 1821 945 1833
rect 974 1821 986 1833
rect 894 1767 906 1779
rect 1015 1821 1027 1833
rect 1154 1841 1166 1853
rect 1134 1821 1146 1833
rect 1074 1781 1086 1793
rect 1254 1841 1266 1853
rect 1175 1821 1187 1833
rect 1234 1821 1246 1833
rect 1275 1821 1287 1833
rect 1414 1801 1426 1813
rect 1374 1781 1386 1793
rect 1534 1841 1546 1853
rect 1514 1821 1526 1833
rect 1493 1801 1505 1813
rect 1435 1767 1447 1779
rect 1473 1767 1485 1779
rect 1555 1821 1567 1833
rect 1614 1781 1626 1793
rect 1794 1841 1806 1853
rect 1773 1821 1785 1833
rect 1714 1767 1726 1779
rect 1814 1821 1826 1833
rect 1834 1801 1846 1813
rect 1874 1787 1886 1799
rect 2021 1858 2033 1870
rect 2003 1824 2015 1836
rect 1954 1781 1966 1793
rect 1974 1782 1986 1794
rect 1875 1750 1887 1762
rect 1994 1768 2006 1780
rect 2055 1858 2067 1870
rect 2035 1838 2047 1850
rect 1997 1736 2009 1748
rect 2019 1736 2031 1748
rect 2083 1844 2095 1856
rect 2107 1844 2119 1856
rect 2067 1740 2079 1752
rect 2135 1812 2147 1824
rect 2121 1773 2133 1785
rect 2194 1801 2206 1813
rect 2234 1801 2246 1813
rect 2314 1801 2326 1813
rect 2254 1781 2266 1793
rect 2373 1821 2385 1833
rect 2334 1767 2346 1779
rect 2414 1801 2426 1813
rect 2454 1801 2466 1813
rect 2494 1801 2506 1813
rect 2534 1801 2546 1813
rect 2574 1801 2586 1813
rect 2633 1821 2645 1833
rect 2594 1767 2606 1779
rect 2694 1787 2706 1799
rect 2774 1801 2786 1813
rect 2814 1801 2826 1813
rect 2834 1801 2846 1813
rect 2734 1787 2746 1799
rect 2893 1821 2905 1833
rect 2854 1767 2866 1779
rect 3121 1844 3133 1856
rect 3173 1858 3185 1870
rect 3145 1844 3157 1856
rect 3014 1801 3026 1813
rect 3054 1801 3066 1813
rect 3093 1812 3105 1824
rect 2934 1781 2946 1793
rect 3107 1773 3119 1785
rect 3161 1740 3173 1752
rect 3207 1858 3219 1870
rect 3193 1838 3205 1850
rect 3225 1824 3237 1836
rect 3254 1782 3266 1794
rect 3314 1801 3326 1813
rect 3234 1768 3246 1780
rect 3209 1736 3221 1748
rect 3231 1736 3243 1748
rect 3274 1781 3286 1793
rect 3373 1821 3385 1833
rect 3334 1767 3346 1779
rect 3414 1787 3426 1799
rect 3541 1844 3553 1856
rect 3593 1858 3605 1870
rect 3565 1844 3577 1856
rect 3513 1812 3525 1824
rect 3454 1787 3466 1799
rect 3527 1773 3539 1785
rect 3581 1740 3593 1752
rect 3627 1858 3639 1870
rect 3613 1838 3625 1850
rect 3645 1824 3657 1836
rect 3674 1782 3686 1794
rect 3763 1818 3775 1830
rect 3734 1801 3746 1813
rect 3654 1768 3666 1780
rect 3629 1736 3641 1748
rect 3651 1736 3663 1748
rect 3694 1781 3706 1793
rect 3834 1787 3846 1799
rect 3915 1821 3927 1833
rect 3874 1787 3886 1799
rect 3763 1750 3775 1762
rect 4015 1821 4027 1833
rect 3974 1801 3986 1813
rect 3954 1767 3966 1779
rect 4074 1801 4086 1813
rect 4054 1767 4066 1779
rect 4133 1819 4145 1831
rect 4114 1801 4126 1813
rect 4094 1781 4106 1793
rect 4481 1844 4493 1856
rect 4533 1858 4545 1870
rect 4505 1844 4517 1856
rect 4234 1781 4246 1793
rect 4133 1752 4145 1764
rect 4274 1781 4286 1793
rect 4254 1767 4266 1779
rect 4374 1801 4386 1813
rect 4414 1801 4426 1813
rect 4453 1812 4465 1824
rect 4294 1767 4306 1779
rect 4467 1773 4479 1785
rect 4521 1740 4533 1752
rect 4567 1858 4579 1870
rect 4553 1838 4565 1850
rect 4585 1824 4597 1836
rect 4614 1782 4626 1794
rect 4594 1768 4606 1780
rect 4569 1736 4581 1748
rect 4591 1736 4603 1748
rect 4634 1781 4646 1793
rect 4694 1787 4706 1799
rect 4734 1787 4746 1799
rect 114 1601 126 1613
rect 54 1587 66 1599
rect 154 1601 166 1613
rect 134 1587 146 1599
rect 174 1547 186 1559
rect 274 1581 286 1593
rect 215 1547 227 1559
rect 194 1527 206 1539
rect 314 1581 326 1593
rect 414 1601 426 1613
rect 375 1547 387 1559
rect 485 1618 497 1630
rect 574 1587 586 1599
rect 434 1567 446 1579
rect 514 1567 526 1579
rect 485 1550 497 1562
rect 594 1547 606 1559
rect 694 1601 706 1613
rect 734 1601 746 1613
rect 714 1587 726 1599
rect 635 1547 647 1559
rect 614 1527 626 1539
rect 794 1547 806 1559
rect 894 1601 906 1613
rect 934 1601 946 1613
rect 914 1587 926 1599
rect 835 1547 847 1559
rect 814 1527 826 1539
rect 994 1547 1006 1559
rect 1154 1601 1166 1613
rect 1035 1547 1047 1559
rect 1115 1547 1127 1559
rect 1014 1527 1026 1539
rect 1174 1567 1186 1579
rect 1194 1547 1206 1559
rect 1294 1601 1306 1613
rect 1334 1601 1346 1613
rect 1314 1587 1326 1599
rect 1235 1547 1247 1559
rect 1214 1527 1226 1539
rect 1434 1587 1446 1599
rect 1454 1547 1466 1559
rect 1554 1601 1566 1613
rect 1594 1601 1606 1613
rect 1574 1587 1586 1599
rect 1495 1547 1507 1559
rect 1474 1527 1486 1539
rect 1654 1547 1666 1559
rect 1774 1601 1786 1613
rect 1754 1567 1766 1579
rect 1695 1547 1707 1559
rect 1674 1527 1686 1539
rect 1894 1601 1906 1613
rect 1813 1547 1825 1559
rect 1934 1601 1946 1613
rect 1914 1587 1926 1599
rect 1954 1587 1966 1599
rect 2014 1547 2026 1559
rect 2174 1601 2186 1613
rect 2055 1547 2067 1559
rect 2135 1547 2147 1559
rect 2034 1527 2046 1539
rect 2214 1587 2226 1599
rect 2194 1567 2206 1579
rect 2307 1595 2319 1607
rect 2293 1556 2305 1568
rect 2361 1628 2373 1640
rect 2321 1524 2333 1536
rect 2345 1524 2357 1536
rect 2409 1632 2421 1644
rect 2431 1632 2443 1644
rect 2393 1530 2405 1542
rect 2373 1510 2385 1522
rect 2434 1600 2446 1612
rect 2454 1586 2466 1598
rect 2474 1587 2486 1599
rect 2425 1544 2437 1556
rect 2407 1510 2419 1522
rect 2574 1601 2586 1613
rect 2535 1547 2547 1559
rect 2653 1618 2665 1630
rect 2594 1567 2606 1579
rect 2654 1581 2666 1593
rect 2794 1601 2806 1613
rect 2694 1567 2706 1579
rect 2714 1567 2726 1579
rect 2754 1567 2766 1579
rect 2834 1601 2846 1613
rect 2814 1587 2826 1599
rect 3014 1587 3026 1599
rect 3074 1587 3086 1599
rect 2914 1567 2926 1579
rect 2954 1567 2966 1579
rect 3114 1601 3126 1613
rect 3094 1567 3106 1579
rect 3194 1581 3206 1593
rect 3153 1547 3165 1559
rect 3234 1581 3246 1593
rect 3294 1581 3306 1593
rect 3334 1581 3346 1593
rect 3414 1601 3426 1613
rect 3375 1547 3387 1559
rect 3474 1587 3486 1599
rect 3517 1632 3529 1644
rect 3539 1632 3551 1644
rect 3514 1600 3526 1612
rect 3434 1567 3446 1579
rect 3494 1586 3506 1598
rect 3523 1544 3535 1556
rect 3555 1530 3567 1542
rect 3541 1510 3553 1522
rect 3587 1628 3599 1640
rect 3641 1595 3653 1607
rect 3694 1587 3706 1599
rect 3655 1556 3667 1568
rect 3603 1524 3615 1536
rect 3575 1510 3587 1522
rect 3627 1524 3639 1536
rect 3794 1587 3806 1599
rect 3874 1601 3886 1613
rect 3835 1547 3847 1559
rect 4134 1601 4146 1613
rect 4074 1587 4086 1599
rect 3894 1567 3906 1579
rect 3914 1567 3926 1579
rect 3954 1567 3966 1579
rect 3994 1567 4006 1579
rect 4034 1567 4046 1579
rect 4174 1601 4186 1613
rect 4154 1587 4166 1599
rect 4314 1601 4326 1613
rect 4234 1567 4246 1579
rect 4274 1567 4286 1579
rect 4354 1601 4366 1613
rect 4334 1587 4346 1599
rect 4414 1587 4426 1599
rect 4474 1587 4486 1599
rect 4574 1587 4586 1599
rect 4614 1601 4626 1613
rect 4594 1567 4606 1579
rect 4694 1581 4706 1593
rect 4653 1547 4665 1559
rect 4734 1581 4746 1593
rect 134 1361 146 1373
rect 114 1341 126 1353
rect 74 1301 86 1313
rect 54 1287 66 1299
rect 94 1287 106 1299
rect 234 1361 246 1373
rect 155 1341 167 1353
rect 214 1341 226 1353
rect 255 1341 267 1353
rect 334 1307 346 1319
rect 394 1321 406 1333
rect 374 1307 386 1319
rect 453 1341 465 1353
rect 414 1287 426 1299
rect 514 1301 526 1313
rect 494 1287 506 1299
rect 594 1321 606 1333
rect 534 1287 546 1299
rect 653 1341 665 1353
rect 614 1287 626 1299
rect 694 1321 706 1333
rect 753 1341 765 1353
rect 714 1287 726 1299
rect 794 1321 806 1333
rect 834 1307 846 1319
rect 914 1307 926 1319
rect 954 1307 966 1319
rect 974 1307 986 1319
rect 835 1270 847 1282
rect 1114 1361 1126 1373
rect 1093 1341 1105 1353
rect 1014 1307 1026 1319
rect 1134 1341 1146 1353
rect 1194 1301 1206 1313
rect 1294 1321 1306 1333
rect 1314 1321 1326 1333
rect 1254 1307 1266 1319
rect 1253 1270 1265 1282
rect 1373 1341 1385 1353
rect 1435 1341 1447 1353
rect 1334 1287 1346 1299
rect 1494 1321 1506 1333
rect 1474 1287 1486 1299
rect 1514 1307 1526 1319
rect 1594 1321 1606 1333
rect 1554 1307 1566 1319
rect 1653 1341 1665 1353
rect 1614 1287 1626 1299
rect 1694 1307 1706 1319
rect 1734 1307 1746 1319
rect 1794 1301 1806 1313
rect 1774 1287 1786 1299
rect 1894 1361 1906 1373
rect 1874 1341 1886 1353
rect 1814 1287 1826 1299
rect 1915 1341 1927 1353
rect 1974 1321 1986 1333
rect 2033 1341 2045 1353
rect 1994 1287 2006 1299
rect 2154 1361 2166 1373
rect 2134 1341 2146 1353
rect 2074 1301 2086 1313
rect 2175 1341 2187 1353
rect 2234 1307 2246 1319
rect 2274 1307 2286 1319
rect 2353 1339 2365 1351
rect 2334 1321 2346 1333
rect 2314 1301 2326 1313
rect 2434 1307 2446 1319
rect 2474 1307 2486 1319
rect 2585 1338 2597 1350
rect 2494 1301 2506 1313
rect 2353 1272 2365 1284
rect 2614 1321 2626 1333
rect 2634 1321 2646 1333
rect 2585 1270 2597 1282
rect 2693 1341 2705 1353
rect 2654 1287 2666 1299
rect 2755 1321 2767 1333
rect 2834 1321 2846 1333
rect 2778 1287 2790 1299
rect 2814 1287 2826 1299
rect 2941 1378 2953 1390
rect 2923 1344 2935 1356
rect 2874 1301 2886 1313
rect 2894 1302 2906 1314
rect 2914 1288 2926 1300
rect 2975 1378 2987 1390
rect 2955 1358 2967 1370
rect 2917 1256 2929 1268
rect 2939 1256 2951 1268
rect 3003 1364 3015 1376
rect 3027 1364 3039 1376
rect 2987 1260 2999 1272
rect 3055 1332 3067 1344
rect 3041 1293 3053 1305
rect 3114 1321 3126 1333
rect 3154 1321 3166 1333
rect 3234 1301 3246 1313
rect 3214 1287 3226 1299
rect 3361 1378 3373 1390
rect 3343 1344 3355 1356
rect 3294 1301 3306 1313
rect 3314 1302 3326 1314
rect 3254 1287 3266 1299
rect 3334 1288 3346 1300
rect 3395 1378 3407 1390
rect 3375 1358 3387 1370
rect 3337 1256 3349 1268
rect 3359 1256 3371 1268
rect 3423 1364 3435 1376
rect 3447 1364 3459 1376
rect 3407 1260 3419 1272
rect 3475 1332 3487 1344
rect 3461 1293 3473 1305
rect 3594 1321 3606 1333
rect 3634 1321 3646 1333
rect 3674 1321 3686 1333
rect 3714 1321 3726 1333
rect 3554 1301 3566 1313
rect 3841 1364 3853 1376
rect 3893 1378 3905 1390
rect 3865 1364 3877 1376
rect 3734 1301 3746 1313
rect 3813 1332 3825 1344
rect 3827 1293 3839 1305
rect 3881 1260 3893 1272
rect 3927 1378 3939 1390
rect 3913 1358 3925 1370
rect 3945 1344 3957 1356
rect 3974 1302 3986 1314
rect 4034 1321 4046 1333
rect 3954 1288 3966 1300
rect 3929 1256 3941 1268
rect 3951 1256 3963 1268
rect 3994 1301 4006 1313
rect 4093 1341 4105 1353
rect 4054 1287 4066 1299
rect 4134 1307 4146 1319
rect 4245 1338 4257 1350
rect 4274 1321 4286 1333
rect 4174 1307 4186 1319
rect 4245 1270 4257 1282
rect 4314 1307 4326 1319
rect 4395 1341 4407 1353
rect 4354 1307 4366 1319
rect 4495 1341 4507 1353
rect 4454 1321 4466 1333
rect 4434 1287 4446 1299
rect 4554 1321 4566 1333
rect 4574 1321 4586 1333
rect 4614 1321 4626 1333
rect 4534 1287 4546 1299
rect 4654 1301 4666 1313
rect 4754 1301 4766 1313
rect 74 1121 86 1133
rect 35 1067 47 1079
rect 134 1121 146 1133
rect 94 1087 106 1099
rect 114 1087 126 1099
rect 173 1067 185 1079
rect 214 1067 226 1079
rect 314 1121 326 1133
rect 354 1121 366 1133
rect 334 1107 346 1119
rect 255 1067 267 1079
rect 234 1047 246 1059
rect 414 1067 426 1079
rect 514 1121 526 1133
rect 554 1121 566 1133
rect 534 1107 546 1119
rect 455 1067 467 1079
rect 434 1047 446 1059
rect 733 1138 745 1150
rect 634 1101 646 1113
rect 674 1101 686 1113
rect 734 1101 746 1113
rect 774 1087 786 1099
rect 833 1067 845 1079
rect 954 1121 966 1133
rect 874 1067 886 1079
rect 915 1067 927 1079
rect 854 1047 866 1059
rect 1014 1121 1026 1133
rect 974 1087 986 1099
rect 994 1087 1006 1099
rect 1154 1121 1166 1133
rect 1053 1067 1065 1079
rect 1115 1067 1127 1079
rect 1313 1138 1325 1150
rect 1214 1101 1226 1113
rect 1174 1087 1186 1099
rect 1254 1101 1266 1113
rect 1314 1101 1326 1113
rect 1374 1101 1386 1113
rect 1354 1087 1366 1099
rect 1494 1121 1506 1133
rect 1414 1101 1426 1113
rect 1534 1101 1546 1113
rect 1574 1101 1586 1113
rect 1614 1101 1626 1113
rect 1654 1101 1666 1113
rect 1674 1067 1686 1079
rect 1794 1101 1806 1113
rect 1715 1067 1727 1079
rect 1694 1047 1706 1059
rect 1834 1101 1846 1113
rect 1854 1067 1866 1079
rect 1954 1101 1966 1113
rect 1895 1067 1907 1079
rect 1874 1047 1886 1059
rect 1994 1101 2006 1113
rect 2075 1121 2087 1133
rect 2113 1121 2125 1133
rect 2054 1087 2066 1099
rect 2133 1087 2145 1099
rect 2193 1067 2205 1079
rect 2274 1101 2286 1113
rect 2234 1067 2246 1079
rect 2214 1047 2226 1059
rect 2334 1121 2346 1133
rect 2314 1101 2326 1113
rect 2374 1121 2386 1133
rect 2354 1107 2366 1119
rect 2474 1107 2486 1119
rect 2514 1101 2526 1113
rect 2554 1101 2566 1113
rect 2618 1121 2630 1133
rect 2654 1121 2666 1133
rect 2595 1087 2607 1099
rect 2723 1138 2735 1150
rect 2794 1107 2806 1119
rect 2837 1152 2849 1164
rect 2859 1152 2871 1164
rect 2834 1120 2846 1132
rect 2674 1087 2686 1099
rect 2694 1087 2706 1099
rect 2723 1070 2735 1082
rect 2814 1106 2826 1118
rect 2843 1064 2855 1076
rect 2875 1050 2887 1062
rect 2861 1030 2873 1042
rect 2907 1148 2919 1160
rect 2961 1115 2973 1127
rect 3014 1101 3026 1113
rect 2975 1076 2987 1088
rect 2923 1044 2935 1056
rect 2895 1030 2907 1042
rect 2947 1044 2959 1056
rect 3054 1101 3066 1113
rect 3154 1121 3166 1133
rect 3115 1067 3127 1079
rect 3345 1138 3357 1150
rect 3423 1138 3435 1150
rect 3174 1087 3186 1099
rect 3214 1087 3226 1099
rect 3374 1087 3386 1099
rect 3394 1087 3406 1099
rect 3345 1070 3357 1082
rect 3494 1121 3506 1133
rect 3530 1124 3542 1136
rect 3570 1124 3582 1136
rect 3610 1124 3622 1136
rect 3423 1070 3435 1082
rect 3694 1121 3706 1133
rect 3730 1124 3742 1136
rect 3770 1124 3782 1136
rect 3810 1124 3822 1136
rect 3903 1138 3915 1150
rect 3954 1101 3966 1113
rect 3874 1087 3886 1099
rect 3903 1070 3915 1082
rect 3994 1101 4006 1113
rect 4067 1115 4079 1127
rect 4053 1076 4065 1088
rect 4121 1148 4133 1160
rect 4081 1044 4093 1056
rect 4105 1044 4117 1056
rect 4169 1152 4181 1164
rect 4191 1152 4203 1164
rect 4153 1050 4165 1062
rect 4133 1030 4145 1042
rect 4194 1120 4206 1132
rect 4214 1106 4226 1118
rect 4234 1107 4246 1119
rect 4185 1064 4197 1076
rect 4167 1030 4179 1042
rect 4274 1101 4286 1113
rect 4314 1101 4326 1113
rect 4374 1121 4386 1133
rect 4354 1087 4366 1099
rect 4474 1101 4486 1113
rect 4413 1067 4425 1079
rect 4514 1101 4526 1113
rect 4554 1121 4566 1133
rect 4534 1087 4546 1099
rect 4593 1067 4605 1079
rect 4634 1067 4646 1079
rect 4675 1067 4687 1079
rect 4654 1047 4666 1059
rect 34 827 46 839
rect 74 827 86 839
rect 215 861 227 873
rect 174 841 186 853
rect 134 827 146 839
rect 133 790 145 802
rect 274 841 286 853
rect 314 841 326 853
rect 254 807 266 819
rect 445 858 457 870
rect 393 841 405 853
rect 474 841 486 853
rect 335 807 347 819
rect 373 807 385 819
rect 445 790 457 802
rect 494 821 506 833
rect 594 821 606 833
rect 734 881 746 893
rect 714 861 726 873
rect 674 821 686 833
rect 654 807 666 819
rect 694 807 706 819
rect 755 861 767 873
rect 894 841 906 853
rect 854 827 866 839
rect 853 790 865 802
rect 914 827 926 839
rect 1054 881 1066 893
rect 1033 861 1045 873
rect 954 827 966 839
rect 1074 861 1086 873
rect 1094 841 1106 853
rect 1254 881 1266 893
rect 1153 861 1165 873
rect 1233 861 1245 873
rect 1114 807 1126 819
rect 1274 861 1286 873
rect 1354 841 1366 853
rect 1294 821 1306 833
rect 1413 861 1425 873
rect 1374 807 1386 819
rect 1474 827 1486 839
rect 1514 827 1526 839
rect 1534 827 1546 839
rect 1635 861 1647 873
rect 1574 827 1586 839
rect 1694 841 1706 853
rect 1714 841 1726 853
rect 1674 807 1686 819
rect 1754 827 1766 839
rect 1755 790 1767 802
rect 1854 821 1866 833
rect 1894 827 1906 839
rect 1934 827 1946 839
rect 2074 881 2086 893
rect 2053 861 2065 873
rect 1954 821 1966 833
rect 2094 861 2106 873
rect 2174 841 2186 853
rect 2114 821 2126 833
rect 2233 861 2245 873
rect 2194 807 2206 819
rect 2334 821 2346 833
rect 2314 807 2326 819
rect 2454 881 2466 893
rect 2434 861 2446 873
rect 2374 821 2386 833
rect 2354 807 2366 819
rect 2475 861 2487 873
rect 2594 881 2606 893
rect 2573 861 2585 873
rect 2614 861 2626 873
rect 2654 821 2666 833
rect 2634 807 2646 819
rect 2754 827 2766 839
rect 2674 807 2686 819
rect 2835 841 2847 853
rect 2794 827 2806 839
rect 2914 841 2926 853
rect 2858 807 2870 819
rect 2894 807 2906 819
rect 3014 841 3026 853
rect 3054 841 3066 853
rect 3094 841 3106 853
rect 3134 841 3146 853
rect 2974 821 2986 833
rect 3214 841 3226 853
rect 3154 821 3166 833
rect 3273 861 3285 873
rect 3234 807 3246 819
rect 3314 827 3326 839
rect 3441 884 3453 896
rect 3493 898 3505 910
rect 3465 884 3477 896
rect 3413 852 3425 864
rect 3354 827 3366 839
rect 3427 813 3439 825
rect 3481 780 3493 792
rect 3527 898 3539 910
rect 3513 878 3525 890
rect 3545 864 3557 876
rect 3574 822 3586 834
rect 3663 858 3675 870
rect 3634 841 3646 853
rect 3554 808 3566 820
rect 3529 776 3541 788
rect 3551 776 3563 788
rect 3594 821 3606 833
rect 3801 898 3813 910
rect 3783 864 3795 876
rect 3734 821 3746 833
rect 3754 822 3766 834
rect 3663 790 3675 802
rect 3774 808 3786 820
rect 3835 898 3847 910
rect 3815 878 3827 890
rect 3777 776 3789 788
rect 3799 776 3811 788
rect 3863 884 3875 896
rect 3887 884 3899 896
rect 3847 780 3859 792
rect 4101 884 4113 896
rect 4153 898 4165 910
rect 4125 884 4137 896
rect 3915 852 3927 864
rect 3975 861 3987 873
rect 3901 813 3913 825
rect 4034 841 4046 853
rect 4073 852 4085 864
rect 4014 807 4026 819
rect 4087 813 4099 825
rect 4141 780 4153 792
rect 4187 898 4199 910
rect 4173 878 4185 890
rect 4205 864 4217 876
rect 4234 822 4246 834
rect 4381 898 4393 910
rect 4363 864 4375 876
rect 4214 808 4226 820
rect 4189 776 4201 788
rect 4211 776 4223 788
rect 4254 821 4266 833
rect 4314 821 4326 833
rect 4334 822 4346 834
rect 4354 808 4366 820
rect 4415 898 4427 910
rect 4395 878 4407 890
rect 4357 776 4369 788
rect 4379 776 4391 788
rect 4443 884 4455 896
rect 4467 884 4479 896
rect 4427 780 4439 792
rect 4495 852 4507 864
rect 4481 813 4493 825
rect 4534 841 4546 853
rect 4593 861 4605 873
rect 4554 807 4566 819
rect 4634 841 4646 853
rect 4693 861 4705 873
rect 4654 807 4666 819
rect 134 641 146 653
rect 34 607 46 619
rect 74 607 86 619
rect 174 641 186 653
rect 154 627 166 639
rect 194 627 206 639
rect 294 641 306 653
rect 334 641 346 653
rect 314 627 326 639
rect 354 587 366 599
rect 514 641 526 653
rect 395 587 407 599
rect 475 587 487 599
rect 374 567 386 579
rect 585 658 597 670
rect 534 607 546 619
rect 614 607 626 619
rect 585 590 597 602
rect 694 641 706 653
rect 655 587 667 599
rect 765 658 777 670
rect 855 658 867 670
rect 854 621 866 633
rect 714 607 726 619
rect 794 607 806 619
rect 814 607 826 619
rect 765 590 777 602
rect 934 641 946 653
rect 914 607 926 619
rect 1074 641 1086 653
rect 973 587 985 599
rect 1035 587 1047 599
rect 1154 641 1166 653
rect 1174 641 1186 653
rect 1094 607 1106 619
rect 1214 641 1226 653
rect 1194 627 1206 639
rect 1314 627 1326 639
rect 1354 641 1366 653
rect 1334 607 1346 619
rect 1454 641 1466 653
rect 1434 607 1446 619
rect 1393 587 1405 599
rect 1574 641 1586 653
rect 1493 587 1505 599
rect 1614 641 1626 653
rect 1634 641 1646 653
rect 1594 627 1606 639
rect 1674 641 1686 653
rect 1654 627 1666 639
rect 1734 587 1746 599
rect 1854 641 1866 653
rect 1834 607 1846 619
rect 1775 587 1787 599
rect 1754 567 1766 579
rect 1974 641 1986 653
rect 1893 587 1905 599
rect 2014 641 2026 653
rect 1994 627 2006 639
rect 2054 641 2066 653
rect 2034 607 2046 619
rect 2093 587 2105 599
rect 2173 587 2185 599
rect 2294 641 2306 653
rect 2214 587 2226 599
rect 2255 587 2267 599
rect 2194 567 2206 579
rect 2354 641 2366 653
rect 2314 607 2326 619
rect 2334 607 2346 619
rect 2393 587 2405 599
rect 2434 587 2446 599
rect 2475 587 2487 599
rect 2534 587 2546 599
rect 2454 567 2466 579
rect 2674 627 2686 639
rect 2575 587 2587 599
rect 2554 567 2566 579
rect 2694 587 2706 599
rect 2814 627 2826 639
rect 2857 672 2869 684
rect 2879 672 2891 684
rect 2854 640 2866 652
rect 2735 587 2747 599
rect 2714 567 2726 579
rect 2834 626 2846 638
rect 2863 584 2875 596
rect 2895 570 2907 582
rect 2881 550 2893 562
rect 2927 668 2939 680
rect 2981 635 2993 647
rect 3054 641 3066 653
rect 2995 596 3007 608
rect 3034 607 3046 619
rect 3134 627 3146 639
rect 3194 627 3206 639
rect 3093 587 3105 599
rect 2943 564 2955 576
rect 2915 550 2927 562
rect 2967 564 2979 576
rect 3254 587 3266 599
rect 3394 627 3406 639
rect 3295 587 3307 599
rect 3274 567 3286 579
rect 3434 621 3446 633
rect 3474 621 3486 633
rect 3554 641 3566 653
rect 3515 587 3527 599
rect 3614 627 3626 639
rect 3657 672 3669 684
rect 3679 672 3691 684
rect 3654 640 3666 652
rect 3574 607 3586 619
rect 3634 626 3646 638
rect 3663 584 3675 596
rect 3695 570 3707 582
rect 3681 550 3693 562
rect 3727 668 3739 680
rect 3781 635 3793 647
rect 3854 641 3866 653
rect 3795 596 3807 608
rect 3834 607 3846 619
rect 3954 621 3966 633
rect 3893 587 3905 599
rect 3743 564 3755 576
rect 3715 550 3727 562
rect 3767 564 3779 576
rect 3994 621 4006 633
rect 4047 635 4059 647
rect 4033 596 4045 608
rect 4101 668 4113 680
rect 4061 564 4073 576
rect 4085 564 4097 576
rect 4149 672 4161 684
rect 4171 672 4183 684
rect 4133 570 4145 582
rect 4113 550 4125 562
rect 4174 640 4186 652
rect 4194 626 4206 638
rect 4214 627 4226 639
rect 4165 584 4177 596
rect 4147 550 4159 562
rect 4254 621 4266 633
rect 4294 621 4306 633
rect 4334 621 4346 633
rect 4374 621 4386 633
rect 4474 641 4486 653
rect 4435 587 4447 599
rect 4534 627 4546 639
rect 4577 672 4589 684
rect 4599 672 4611 684
rect 4574 640 4586 652
rect 4494 607 4506 619
rect 4554 626 4566 638
rect 4583 584 4595 596
rect 4615 570 4627 582
rect 4601 550 4613 562
rect 4647 668 4659 680
rect 4701 635 4713 647
rect 4715 596 4727 608
rect 4663 564 4675 576
rect 4635 550 4647 562
rect 4687 564 4699 576
rect 14 347 26 359
rect 54 347 66 359
rect 94 347 106 359
rect 134 347 146 359
rect 194 347 206 359
rect 234 347 246 359
rect 274 347 286 359
rect 314 347 326 359
rect 414 361 426 373
rect 374 347 386 359
rect 373 310 385 322
rect 454 347 466 359
rect 574 401 586 413
rect 553 381 565 393
rect 494 347 506 359
rect 594 381 606 393
rect 634 361 646 373
rect 713 361 725 373
rect 754 361 766 373
rect 794 361 806 373
rect 655 327 667 339
rect 693 327 705 339
rect 834 347 846 359
rect 874 347 886 359
rect 894 347 906 359
rect 934 347 946 359
rect 994 347 1006 359
rect 1034 347 1046 359
rect 1074 347 1086 359
rect 1154 361 1166 373
rect 1114 347 1126 359
rect 1233 361 1245 373
rect 1254 361 1266 373
rect 1175 327 1187 339
rect 1213 327 1225 339
rect 1313 381 1325 393
rect 1274 327 1286 339
rect 1374 361 1386 373
rect 1414 361 1426 373
rect 1434 361 1446 373
rect 1493 381 1505 393
rect 1454 327 1466 339
rect 1534 341 1546 353
rect 1654 341 1666 353
rect 1634 327 1646 339
rect 1774 401 1786 413
rect 1754 381 1766 393
rect 1694 341 1706 353
rect 1674 327 1686 339
rect 1795 381 1807 393
rect 1874 341 1886 353
rect 1854 327 1866 339
rect 1954 347 1966 359
rect 1894 327 1906 339
rect 1994 347 2006 359
rect 2034 347 2046 359
rect 2074 347 2086 359
rect 2114 347 2126 359
rect 2214 361 2226 373
rect 2254 361 2266 373
rect 2154 347 2166 359
rect 2294 347 2306 359
rect 2354 361 2366 373
rect 2454 401 2466 413
rect 2434 381 2446 393
rect 2394 361 2406 373
rect 2334 347 2346 359
rect 2475 381 2487 393
rect 2654 401 2666 413
rect 2633 381 2645 393
rect 2574 341 2586 353
rect 2674 381 2686 393
rect 2714 341 2726 353
rect 2694 327 2706 339
rect 2794 361 2806 373
rect 2834 361 2846 373
rect 2734 327 2746 339
rect 2894 347 2906 359
rect 2975 381 2987 393
rect 2934 347 2946 359
rect 3075 381 3087 393
rect 3034 361 3046 373
rect 3014 327 3026 339
rect 3134 361 3146 373
rect 3174 361 3186 373
rect 3214 361 3226 373
rect 3114 327 3126 339
rect 3315 381 3327 393
rect 3274 341 3286 353
rect 3374 361 3386 373
rect 3354 327 3366 339
rect 3454 341 3466 353
rect 3434 327 3446 339
rect 3514 361 3526 373
rect 3554 361 3566 373
rect 3474 327 3486 339
rect 3613 379 3625 391
rect 3594 361 3606 373
rect 3574 341 3586 353
rect 3674 347 3686 359
rect 3714 347 3726 359
rect 3754 347 3766 359
rect 3613 312 3625 324
rect 3855 381 3867 393
rect 3794 347 3806 359
rect 3914 361 3926 373
rect 3894 327 3906 339
rect 4101 404 4113 416
rect 4153 418 4165 430
rect 4125 404 4137 416
rect 4073 372 4085 384
rect 3974 341 3986 353
rect 4034 341 4046 353
rect 4087 333 4099 345
rect 4141 300 4153 312
rect 4187 418 4199 430
rect 4173 398 4185 410
rect 4205 384 4217 396
rect 4234 342 4246 354
rect 4214 328 4226 340
rect 4189 296 4201 308
rect 4211 296 4223 308
rect 4254 341 4266 353
rect 4314 347 4326 359
rect 4395 381 4407 393
rect 4354 347 4366 359
rect 4454 361 4466 373
rect 4434 327 4446 339
rect 4581 404 4593 416
rect 4633 418 4645 430
rect 4605 404 4617 416
rect 4553 372 4565 384
rect 4514 341 4526 353
rect 4567 333 4579 345
rect 4621 300 4633 312
rect 4667 418 4679 430
rect 4653 398 4665 410
rect 4685 384 4697 396
rect 4714 342 4726 354
rect 4694 328 4706 340
rect 4669 296 4681 308
rect 4691 296 4703 308
rect 4734 341 4746 353
rect 53 107 65 119
rect 114 161 126 173
rect 154 161 166 173
rect 134 147 146 159
rect 94 107 106 119
rect 74 87 86 99
rect 274 161 286 173
rect 235 107 247 119
rect 334 161 346 173
rect 294 127 306 139
rect 314 127 326 139
rect 373 107 385 119
rect 453 107 465 119
rect 494 107 506 119
rect 514 107 526 119
rect 474 87 486 99
rect 614 161 626 173
rect 654 161 666 173
rect 634 147 646 159
rect 555 107 567 119
rect 534 87 546 99
rect 754 161 766 173
rect 794 161 806 173
rect 774 147 786 159
rect 814 147 826 159
rect 934 161 946 173
rect 895 107 907 119
rect 1014 147 1026 159
rect 954 127 966 139
rect 1054 161 1066 173
rect 1034 127 1046 139
rect 1154 161 1166 173
rect 1134 127 1146 139
rect 1093 107 1105 119
rect 1193 107 1205 119
rect 1234 107 1246 119
rect 1275 107 1287 119
rect 1334 107 1346 119
rect 1254 87 1266 99
rect 1474 161 1486 173
rect 1375 107 1387 119
rect 1354 87 1366 99
rect 1514 161 1526 173
rect 1494 147 1506 159
rect 1534 107 1546 119
rect 1674 161 1686 173
rect 1575 107 1587 119
rect 1554 87 1566 99
rect 1714 161 1726 173
rect 1694 147 1706 159
rect 1734 107 1746 119
rect 1834 141 1846 153
rect 1775 107 1787 119
rect 1754 87 1766 99
rect 1874 141 1886 153
rect 1943 178 1955 190
rect 2033 178 2045 190
rect 1914 127 1926 139
rect 1943 110 1955 122
rect 2034 141 2046 153
rect 2123 178 2135 190
rect 2074 127 2086 139
rect 2094 127 2106 139
rect 2123 110 2135 122
rect 2174 107 2186 119
rect 2295 161 2307 173
rect 2333 161 2345 173
rect 2275 127 2287 139
rect 2215 107 2227 119
rect 2194 87 2206 99
rect 2414 161 2426 173
rect 2354 127 2366 139
rect 2394 127 2406 139
rect 2534 161 2546 173
rect 2453 107 2465 119
rect 2574 161 2586 173
rect 2554 147 2566 159
rect 2614 161 2626 173
rect 2594 127 2606 139
rect 2694 147 2706 159
rect 2653 107 2665 119
rect 2754 107 2766 119
rect 2854 147 2866 159
rect 2934 147 2946 159
rect 2977 192 2989 204
rect 2999 192 3011 204
rect 2974 160 2986 172
rect 2795 107 2807 119
rect 2774 87 2786 99
rect 2954 146 2966 158
rect 2983 104 2995 116
rect 3015 90 3027 102
rect 3001 70 3013 82
rect 3047 188 3059 200
rect 3101 155 3113 167
rect 3154 147 3166 159
rect 3115 116 3127 128
rect 3063 84 3075 96
rect 3035 70 3047 82
rect 3087 84 3099 96
rect 3254 147 3266 159
rect 3294 147 3306 159
rect 3337 192 3349 204
rect 3359 192 3371 204
rect 3334 160 3346 172
rect 3314 146 3326 158
rect 3343 104 3355 116
rect 3375 90 3387 102
rect 3361 70 3373 82
rect 3407 188 3419 200
rect 3461 155 3473 167
rect 3475 116 3487 128
rect 3534 127 3546 139
rect 3574 127 3586 139
rect 3627 155 3639 167
rect 3613 116 3625 128
rect 3423 84 3435 96
rect 3395 70 3407 82
rect 3447 84 3459 96
rect 3681 188 3693 200
rect 3641 84 3653 96
rect 3665 84 3677 96
rect 3729 192 3741 204
rect 3751 192 3763 204
rect 3713 90 3725 102
rect 3693 70 3705 82
rect 3754 160 3766 172
rect 3774 146 3786 158
rect 3794 147 3806 159
rect 3834 147 3846 159
rect 3745 104 3757 116
rect 3727 70 3739 82
rect 3914 161 3926 173
rect 3894 127 3906 139
rect 4254 161 4266 173
rect 3994 127 4006 139
rect 3953 107 3965 119
rect 4034 127 4046 139
rect 4074 127 4086 139
rect 4114 127 4126 139
rect 4174 127 4186 139
rect 4214 127 4226 139
rect 4234 127 4246 139
rect 4354 141 4366 153
rect 4293 107 4305 119
rect 4394 141 4406 153
rect 4454 147 4466 159
rect 4554 141 4566 153
rect 4474 127 4486 139
rect 4514 127 4526 139
rect 4594 141 4606 153
rect 4674 147 4686 159
rect 4694 141 4706 153
rect 4734 141 4746 153
<< metal1 >>
rect -62 4338 -2 4578
rect 4 4576 4842 4578
rect 4776 4564 4842 4576
rect 4 4562 4842 4564
rect 38 4556 50 4562
rect 88 4556 100 4562
rect 190 4556 202 4562
rect 34 4516 60 4527
rect 34 4473 42 4516
rect 136 4498 154 4500
rect 136 4489 166 4498
rect 218 4556 230 4562
rect 390 4556 402 4562
rect 266 4498 284 4500
rect 254 4489 284 4498
rect 136 4461 144 4489
rect 276 4461 284 4489
rect 336 4498 354 4500
rect 336 4489 366 4498
rect 420 4556 432 4562
rect 470 4556 482 4562
rect 537 4556 549 4562
rect 637 4556 649 4562
rect 790 4556 802 4562
rect 460 4516 486 4527
rect 336 4461 344 4489
rect 478 4473 486 4516
rect 529 4516 557 4522
rect 517 4513 569 4516
rect 629 4516 657 4522
rect 577 4502 585 4516
rect 617 4513 669 4516
rect 677 4502 685 4516
rect 560 4495 585 4502
rect 660 4495 685 4502
rect 736 4498 754 4500
rect 34 4424 42 4459
rect 63 4418 103 4424
rect 91 4416 103 4418
rect 135 4392 142 4447
rect 278 4392 285 4447
rect 135 4386 182 4392
rect 135 4384 143 4386
rect 171 4384 182 4386
rect 238 4386 285 4392
rect 238 4384 249 4386
rect 71 4338 83 4344
rect 151 4338 163 4344
rect 191 4338 203 4344
rect 277 4384 285 4386
rect 335 4392 342 4447
rect 478 4424 486 4459
rect 497 4447 503 4493
rect 559 4473 567 4495
rect 659 4473 667 4495
rect 736 4489 766 4498
rect 818 4556 830 4562
rect 919 4556 931 4562
rect 998 4556 1010 4562
rect 1100 4556 1112 4562
rect 1150 4556 1162 4562
rect 1249 4556 1261 4562
rect 949 4508 961 4516
rect 937 4502 961 4508
rect 866 4498 884 4500
rect 854 4489 884 4498
rect 736 4461 744 4489
rect 876 4461 884 4489
rect 553 4424 561 4459
rect 653 4424 661 4459
rect 417 4418 457 4424
rect 417 4416 429 4418
rect 335 4386 382 4392
rect 335 4384 343 4386
rect 371 4384 382 4386
rect 217 4338 229 4344
rect 257 4338 269 4344
rect 351 4338 363 4344
rect 391 4338 403 4344
rect 437 4338 449 4344
rect 522 4338 534 4344
rect 572 4338 584 4344
rect 735 4392 742 4447
rect 937 4453 945 4502
rect 1140 4516 1166 4527
rect 1046 4498 1064 4500
rect 1034 4489 1064 4498
rect 1056 4461 1064 4489
rect 1158 4473 1166 4516
rect 1291 4556 1303 4562
rect 1331 4556 1343 4562
rect 1411 4556 1423 4562
rect 1509 4556 1521 4562
rect 1219 4508 1231 4516
rect 1219 4502 1243 4508
rect 878 4392 885 4447
rect 735 4386 782 4392
rect 735 4384 743 4386
rect 771 4384 782 4386
rect 838 4386 885 4392
rect 838 4384 849 4386
rect 622 4338 634 4344
rect 672 4338 684 4344
rect 751 4338 763 4344
rect 791 4338 803 4344
rect 877 4384 885 4386
rect 937 4384 945 4439
rect 1058 4392 1065 4447
rect 1158 4424 1166 4459
rect 1235 4453 1243 4502
rect 1313 4493 1320 4536
rect 1375 4502 1383 4516
rect 1403 4516 1431 4522
rect 1391 4513 1443 4516
rect 1537 4556 1549 4562
rect 1577 4556 1589 4562
rect 1618 4556 1630 4562
rect 1738 4556 1750 4562
rect 1788 4556 1800 4562
rect 1479 4508 1491 4516
rect 1479 4502 1503 4508
rect 1375 4495 1400 4502
rect 1018 4386 1065 4392
rect 1018 4384 1029 4386
rect 817 4338 829 4344
rect 857 4338 869 4344
rect 917 4338 929 4344
rect 957 4338 969 4344
rect 1057 4384 1065 4386
rect 1097 4418 1137 4424
rect 1097 4416 1109 4418
rect 1235 4384 1243 4439
rect 1313 4431 1320 4479
rect 1393 4473 1401 4495
rect 1303 4424 1320 4431
rect 1399 4424 1407 4459
rect 1495 4453 1503 4502
rect 1560 4493 1567 4536
rect 1734 4516 1760 4527
rect 1817 4556 1829 4562
rect 1911 4556 1923 4562
rect 1940 4556 1952 4562
rect 1990 4556 2002 4562
rect 1666 4498 1684 4500
rect 1654 4489 1684 4498
rect 997 4338 1009 4344
rect 1037 4338 1049 4344
rect 1117 4338 1129 4344
rect 1211 4338 1223 4344
rect 1251 4338 1263 4344
rect 1331 4338 1343 4344
rect 1495 4384 1503 4439
rect 1560 4431 1567 4479
rect 1676 4461 1684 4489
rect 1734 4473 1742 4516
rect 1836 4481 1844 4536
rect 1896 4481 1904 4536
rect 2037 4556 2049 4562
rect 2077 4556 2089 4562
rect 2117 4556 2129 4562
rect 2197 4556 2209 4562
rect 2351 4556 2363 4562
rect 2397 4556 2405 4562
rect 2437 4556 2449 4562
rect 2500 4556 2512 4562
rect 2550 4556 2562 4562
rect 1980 4516 2006 4527
rect 1998 4473 2006 4516
rect 2060 4493 2067 4536
rect 2136 4481 2144 4536
rect 2189 4516 2217 4522
rect 2177 4513 2229 4516
rect 2303 4550 2331 4556
rect 2343 4516 2371 4520
rect 2237 4502 2245 4516
rect 2220 4495 2245 4502
rect 2315 4506 2321 4516
rect 2331 4514 2383 4516
rect 2423 4508 2429 4536
rect 2632 4556 2644 4562
rect 2688 4556 2700 4562
rect 2741 4556 2753 4562
rect 2803 4556 2815 4562
rect 2851 4556 2863 4562
rect 2909 4556 2921 4562
rect 2991 4556 3003 4562
rect 3071 4556 3083 4562
rect 3131 4556 3143 4562
rect 3171 4556 3183 4562
rect 3251 4556 3263 4562
rect 3311 4556 3323 4562
rect 3351 4556 3363 4562
rect 3411 4556 3423 4562
rect 3459 4556 3471 4562
rect 3517 4556 3529 4562
rect 3565 4556 3577 4562
rect 3627 4556 3639 4562
rect 3697 4556 3709 4562
rect 3779 4556 3791 4562
rect 3871 4556 3883 4562
rect 3911 4556 3923 4562
rect 3951 4556 3963 4562
rect 3991 4556 4003 4562
rect 4031 4556 4043 4562
rect 4089 4556 4101 4562
rect 4139 4556 4151 4562
rect 4217 4556 4229 4562
rect 4297 4556 4309 4562
rect 4399 4556 4411 4562
rect 4457 4556 4469 4562
rect 4505 4556 4517 4562
rect 4567 4556 4579 4562
rect 4639 4556 4651 4562
rect 4699 4556 4711 4562
rect 2540 4516 2566 4527
rect 2760 4536 2773 4542
rect 2760 4530 2767 4536
rect 2825 4524 2832 4536
rect 2315 4499 2344 4506
rect 2423 4502 2433 4508
rect 1560 4424 1577 4431
rect 1376 4338 1388 4344
rect 1426 4338 1438 4344
rect 1471 4338 1483 4344
rect 1511 4338 1523 4344
rect 1678 4392 1685 4447
rect 1734 4424 1742 4459
rect 1638 4386 1685 4392
rect 1638 4384 1649 4386
rect 1677 4384 1685 4386
rect 1763 4418 1803 4424
rect 1791 4416 1803 4418
rect 1836 4384 1844 4467
rect 1896 4384 1904 4467
rect 1998 4424 2006 4459
rect 2060 4431 2067 4479
rect 2060 4424 2077 4431
rect 1937 4418 1977 4424
rect 1937 4416 1949 4418
rect 2136 4384 2144 4467
rect 2219 4473 2227 4495
rect 2336 4473 2344 4499
rect 2213 4424 2221 4459
rect 2335 4424 2343 4459
rect 2438 4441 2444 4496
rect 2460 4481 2467 4516
rect 2558 4473 2566 4516
rect 2397 4432 2433 4440
rect 2397 4424 2405 4432
rect 1537 4338 1549 4344
rect 1617 4338 1629 4344
rect 1657 4338 1669 4344
rect 1771 4338 1783 4344
rect 1817 4338 1829 4344
rect 1911 4338 1923 4344
rect 1957 4338 1969 4344
rect 2037 4338 2049 4344
rect 2117 4338 2129 4344
rect 2182 4338 2194 4344
rect 2232 4338 2244 4344
rect 2454 4423 2463 4467
rect 2660 4473 2667 4516
rect 2558 4424 2566 4459
rect 2653 4436 2659 4459
rect 2632 4430 2659 4436
rect 2721 4432 2727 4516
rect 2811 4517 2832 4524
rect 2882 4530 2889 4536
rect 2882 4522 2893 4530
rect 2779 4506 2786 4512
rect 2847 4506 2853 4508
rect 2779 4500 2853 4506
rect 2935 4501 2943 4516
rect 2779 4492 2786 4500
rect 2740 4484 2774 4492
rect 2740 4479 2746 4484
rect 2766 4466 2793 4473
rect 2632 4424 2644 4430
rect 2721 4424 2783 4432
rect 2795 4428 2839 4434
rect 2459 4414 2463 4423
rect 2497 4418 2537 4424
rect 2497 4416 2509 4418
rect 2623 4344 2651 4350
rect 2663 4416 2691 4422
rect 2777 4410 2815 4418
rect 2833 4414 2839 4428
rect 2847 4428 2853 4500
rect 2927 4487 2943 4501
rect 2913 4473 2927 4487
rect 2847 4422 2887 4428
rect 2907 4428 2921 4436
rect 2935 4424 2943 4487
rect 2976 4481 2984 4536
rect 3035 4502 3043 4516
rect 3063 4516 3091 4522
rect 3051 4513 3103 4516
rect 3117 4517 3133 4523
rect 3035 4495 3060 4502
rect 3053 4473 3061 4495
rect 2777 4404 2785 4410
rect 2833 4408 2863 4414
rect 2881 4404 2887 4422
rect 2767 4390 2785 4404
rect 2813 4390 2835 4402
rect 2777 4384 2785 4390
rect 2827 4384 2839 4390
rect 2881 4364 2893 4398
rect 2976 4384 2984 4467
rect 3059 4424 3067 4459
rect 3117 4447 3123 4517
rect 3153 4493 3160 4536
rect 3215 4502 3223 4516
rect 3243 4516 3271 4522
rect 3231 4513 3283 4516
rect 3215 4495 3240 4502
rect 3153 4431 3160 4479
rect 3233 4473 3241 4495
rect 3333 4493 3340 4536
rect 3396 4481 3404 4536
rect 3607 4536 3620 4542
rect 3491 4530 3498 4536
rect 3487 4522 3498 4530
rect 3548 4524 3555 4536
rect 3613 4530 3620 4536
rect 3437 4501 3445 4516
rect 3548 4517 3569 4524
rect 3527 4506 3533 4508
rect 3594 4506 3601 4512
rect 3143 4424 3160 4431
rect 3239 4424 3247 4459
rect 3333 4431 3340 4479
rect 3437 4487 3453 4501
rect 3527 4500 3601 4506
rect 3323 4424 3340 4431
rect 2301 4338 2313 4344
rect 2371 4338 2383 4344
rect 2427 4338 2439 4344
rect 2517 4338 2529 4344
rect 2671 4338 2683 4344
rect 2741 4338 2753 4344
rect 2807 4338 2819 4344
rect 2853 4338 2865 4344
rect 2911 4338 2923 4344
rect 2991 4338 3003 4344
rect 3036 4338 3048 4344
rect 3086 4338 3098 4344
rect 3171 4338 3183 4344
rect 3396 4384 3404 4467
rect 3437 4424 3445 4487
rect 3453 4473 3467 4487
rect 3459 4428 3473 4436
rect 3527 4428 3533 4500
rect 3594 4492 3601 4500
rect 3606 4484 3640 4492
rect 3634 4479 3640 4484
rect 3587 4466 3614 4473
rect 3493 4422 3533 4428
rect 3541 4428 3585 4434
rect 3493 4404 3499 4422
rect 3541 4414 3547 4428
rect 3653 4432 3659 4516
rect 3689 4516 3717 4522
rect 3677 4513 3729 4516
rect 3737 4502 3745 4516
rect 3809 4508 3821 4516
rect 3892 4510 3904 4516
rect 3932 4510 3944 4516
rect 3971 4510 3983 4516
rect 4012 4510 4024 4516
rect 3886 4509 3904 4510
rect 3720 4495 3745 4502
rect 3797 4502 3821 4508
rect 3885 4502 3904 4509
rect 3918 4502 3944 4510
rect 3958 4502 3983 4510
rect 3997 4502 4024 4510
rect 3719 4473 3727 4495
rect 3597 4424 3659 4432
rect 3713 4424 3721 4459
rect 3797 4453 3805 4502
rect 3885 4481 3892 4502
rect 3918 4496 3926 4502
rect 3958 4496 3966 4502
rect 3997 4496 4005 4502
rect 3910 4484 3926 4496
rect 3950 4484 3966 4496
rect 3990 4484 4005 4496
rect 3887 4467 3892 4481
rect 3517 4408 3547 4414
rect 3565 4410 3603 4418
rect 3595 4404 3603 4410
rect 3487 4364 3499 4398
rect 3545 4390 3567 4402
rect 3595 4390 3613 4404
rect 3541 4384 3553 4390
rect 3595 4384 3603 4390
rect 3797 4384 3805 4439
rect 3885 4438 3892 4467
rect 3918 4438 3926 4484
rect 3958 4438 3966 4484
rect 3997 4438 4005 4484
rect 4071 4473 4079 4516
rect 4111 4510 4119 4536
rect 4097 4504 4119 4510
rect 4169 4508 4181 4516
rect 4097 4498 4100 4504
rect 4071 4459 4073 4473
rect 3885 4430 3903 4438
rect 3918 4430 3943 4438
rect 3958 4430 3983 4438
rect 3997 4430 4023 4438
rect 3891 4424 3903 4430
rect 3931 4424 3943 4430
rect 3971 4424 3983 4430
rect 4011 4424 4023 4430
rect 4071 4424 4079 4459
rect 4093 4442 4100 4498
rect 4157 4502 4181 4508
rect 4157 4453 4165 4502
rect 4236 4481 4244 4536
rect 4289 4516 4317 4522
rect 4277 4513 4329 4516
rect 4547 4536 4560 4542
rect 4431 4530 4438 4536
rect 4427 4522 4438 4530
rect 4488 4524 4495 4536
rect 4553 4530 4560 4536
rect 4337 4502 4345 4516
rect 4320 4495 4345 4502
rect 4377 4501 4385 4516
rect 4488 4517 4509 4524
rect 4467 4506 4473 4508
rect 4534 4506 4541 4512
rect 4097 4436 4100 4442
rect 4097 4430 4123 4436
rect 3216 4338 3228 4344
rect 3266 4338 3278 4344
rect 3351 4338 3363 4344
rect 3411 4338 3423 4344
rect 3457 4338 3469 4344
rect 3515 4338 3527 4344
rect 3561 4338 3573 4344
rect 3627 4338 3639 4344
rect 3682 4338 3694 4344
rect 3732 4338 3744 4344
rect 3777 4338 3789 4344
rect 3817 4338 3829 4344
rect 4115 4384 4123 4430
rect 4157 4384 4165 4439
rect 4236 4384 4244 4467
rect 4319 4473 4327 4495
rect 4377 4487 4393 4501
rect 4467 4500 4541 4506
rect 4313 4424 4321 4459
rect 4377 4424 4385 4487
rect 4393 4473 4407 4487
rect 4399 4428 4413 4436
rect 3871 4338 3883 4344
rect 3911 4338 3923 4344
rect 3951 4338 3963 4344
rect 3991 4338 4003 4344
rect 4031 4338 4043 4344
rect 4089 4338 4101 4344
rect 4137 4338 4149 4344
rect 4177 4338 4189 4344
rect 4467 4428 4473 4500
rect 4534 4492 4541 4500
rect 4546 4484 4580 4492
rect 4574 4479 4580 4484
rect 4527 4466 4554 4473
rect 4433 4422 4473 4428
rect 4481 4428 4525 4434
rect 4433 4404 4439 4422
rect 4481 4414 4487 4428
rect 4593 4432 4599 4516
rect 4621 4510 4629 4536
rect 4621 4504 4643 4510
rect 4640 4498 4643 4504
rect 4640 4442 4647 4498
rect 4661 4473 4669 4516
rect 4729 4508 4741 4516
rect 4717 4502 4741 4508
rect 4667 4459 4669 4473
rect 4640 4436 4643 4442
rect 4537 4424 4599 4432
rect 4457 4408 4487 4414
rect 4505 4410 4543 4418
rect 4535 4404 4543 4410
rect 4427 4364 4439 4398
rect 4485 4390 4507 4402
rect 4535 4390 4553 4404
rect 4481 4384 4493 4390
rect 4535 4384 4543 4390
rect 4617 4430 4643 4436
rect 4617 4384 4625 4430
rect 4661 4424 4669 4459
rect 4717 4453 4725 4502
rect 4717 4384 4725 4439
rect 4217 4338 4229 4344
rect 4282 4338 4294 4344
rect 4332 4338 4344 4344
rect 4397 4338 4409 4344
rect 4455 4338 4467 4344
rect 4501 4338 4513 4344
rect 4567 4338 4579 4344
rect 4639 4338 4651 4344
rect 4697 4338 4709 4344
rect 4737 4338 4749 4344
rect -62 4336 4776 4338
rect -62 4324 4 4336
rect -62 4322 4776 4324
rect -62 3858 -2 4322
rect 31 4316 43 4322
rect 71 4316 83 4322
rect 117 4316 129 4322
rect 211 4316 223 4322
rect 251 4316 263 4322
rect 331 4316 343 4322
rect 55 4221 63 4276
rect 97 4242 109 4244
rect 97 4236 137 4242
rect 55 4158 63 4207
rect 158 4201 166 4236
rect 235 4221 243 4276
rect 376 4316 388 4322
rect 426 4316 438 4322
rect 462 4316 474 4322
rect 512 4316 524 4322
rect 591 4316 603 4322
rect 671 4316 683 4322
rect 751 4316 763 4322
rect 303 4229 320 4236
rect 39 4152 63 4158
rect 39 4144 51 4152
rect 158 4144 166 4187
rect 235 4158 243 4207
rect 69 4098 81 4104
rect 140 4133 166 4144
rect 219 4152 243 4158
rect 313 4181 320 4229
rect 399 4201 407 4236
rect 493 4201 501 4236
rect 219 4144 231 4152
rect 313 4124 320 4167
rect 393 4165 401 4187
rect 576 4193 584 4276
rect 777 4316 789 4322
rect 817 4316 829 4322
rect 951 4316 963 4322
rect 1031 4316 1043 4322
rect 1071 4316 1083 4322
rect 691 4242 703 4244
rect 663 4236 703 4242
rect 634 4201 642 4236
rect 499 4165 507 4187
rect 736 4193 744 4276
rect 798 4274 809 4276
rect 837 4274 845 4276
rect 798 4268 845 4274
rect 838 4213 845 4268
rect 903 4310 931 4316
rect 943 4238 971 4244
rect 1015 4274 1023 4276
rect 1097 4316 1109 4322
rect 1137 4316 1149 4322
rect 1211 4316 1223 4322
rect 1251 4316 1263 4322
rect 1311 4316 1323 4322
rect 1351 4316 1363 4322
rect 1051 4274 1062 4276
rect 1015 4268 1062 4274
rect 1118 4274 1129 4276
rect 1157 4274 1165 4276
rect 1118 4268 1165 4274
rect 912 4230 924 4236
rect 912 4224 939 4230
rect 933 4201 939 4224
rect 1015 4213 1022 4268
rect 375 4158 400 4165
rect 500 4158 525 4165
rect 375 4144 383 4158
rect 100 4098 112 4104
rect 150 4098 162 4104
rect 249 4098 261 4104
rect 391 4144 443 4147
rect 403 4138 431 4144
rect 457 4144 509 4147
rect 469 4138 497 4144
rect 517 4144 525 4158
rect 576 4124 584 4179
rect 634 4144 642 4187
rect 634 4133 660 4144
rect 291 4098 303 4104
rect 331 4098 343 4104
rect 411 4098 423 4104
rect 477 4098 489 4104
rect 591 4098 603 4104
rect 736 4124 744 4179
rect 836 4171 844 4199
rect 638 4098 650 4104
rect 688 4098 700 4104
rect 751 4098 763 4104
rect 814 4162 844 4171
rect 826 4160 844 4162
rect 940 4144 947 4187
rect 1158 4213 1165 4268
rect 1235 4221 1243 4276
rect 1295 4274 1303 4276
rect 1391 4316 1403 4322
rect 1431 4316 1443 4322
rect 1457 4316 1469 4322
rect 1497 4316 1509 4322
rect 1611 4316 1623 4322
rect 1691 4316 1703 4322
rect 1331 4274 1342 4276
rect 1295 4268 1342 4274
rect 1295 4213 1302 4268
rect 1415 4221 1423 4276
rect 1478 4274 1489 4276
rect 1517 4274 1525 4276
rect 1478 4268 1525 4274
rect 1016 4171 1024 4199
rect 1156 4171 1164 4199
rect 1016 4162 1046 4171
rect 1016 4160 1034 4162
rect 778 4098 790 4104
rect 912 4098 924 4104
rect 968 4098 980 4104
rect 1070 4098 1082 4104
rect 1134 4162 1164 4171
rect 1146 4160 1164 4162
rect 1235 4158 1243 4207
rect 1296 4171 1304 4199
rect 1296 4162 1326 4171
rect 1296 4160 1314 4162
rect 1219 4152 1243 4158
rect 1219 4144 1231 4152
rect 1415 4158 1423 4207
rect 1518 4213 1525 4268
rect 1722 4316 1734 4322
rect 1772 4316 1784 4322
rect 1831 4316 1843 4322
rect 1871 4316 1883 4322
rect 1897 4316 1909 4322
rect 1957 4316 1969 4322
rect 1997 4316 2009 4322
rect 2057 4316 2069 4322
rect 2097 4316 2109 4322
rect 2181 4316 2193 4322
rect 2247 4316 2259 4322
rect 2293 4316 2305 4322
rect 2351 4316 2363 4322
rect 2419 4316 2431 4322
rect 2511 4316 2523 4322
rect 2591 4316 2603 4322
rect 2637 4316 2649 4322
rect 2695 4316 2707 4322
rect 2741 4316 2753 4322
rect 2807 4316 2819 4322
rect 2857 4316 2869 4322
rect 2971 4316 2983 4322
rect 1583 4229 1600 4236
rect 1663 4229 1680 4236
rect 1516 4171 1524 4199
rect 1399 4152 1423 4158
rect 1399 4144 1411 4152
rect 1098 4098 1110 4104
rect 1249 4098 1261 4104
rect 1350 4098 1362 4104
rect 1429 4098 1441 4104
rect 1494 4162 1524 4171
rect 1506 4160 1524 4162
rect 1593 4181 1600 4229
rect 1673 4181 1680 4229
rect 1753 4201 1761 4236
rect 1855 4221 1863 4276
rect 1593 4124 1600 4167
rect 1673 4124 1680 4167
rect 1759 4165 1767 4187
rect 1760 4158 1785 4165
rect 1855 4158 1863 4207
rect 1916 4193 1924 4276
rect 1978 4274 1989 4276
rect 2017 4274 2025 4276
rect 1978 4268 2025 4274
rect 2078 4274 2089 4276
rect 2117 4274 2125 4276
rect 2078 4268 2125 4274
rect 2018 4213 2025 4268
rect 2118 4213 2125 4268
rect 2217 4270 2225 4276
rect 2267 4270 2279 4276
rect 2207 4256 2225 4270
rect 2253 4258 2275 4270
rect 2321 4262 2333 4296
rect 2217 4250 2225 4256
rect 2217 4242 2255 4250
rect 2273 4246 2303 4252
rect 2161 4228 2223 4236
rect 1717 4144 1769 4147
rect 1458 4098 1470 4104
rect 1571 4098 1583 4104
rect 1611 4098 1623 4104
rect 1729 4138 1757 4144
rect 1777 4144 1785 4158
rect 1839 4152 1863 4158
rect 1839 4144 1851 4152
rect 1916 4124 1924 4179
rect 2016 4171 2024 4199
rect 2116 4171 2124 4199
rect 1651 4098 1663 4104
rect 1691 4098 1703 4104
rect 1737 4098 1749 4104
rect 1869 4098 1881 4104
rect 1994 4162 2024 4171
rect 2006 4160 2024 4162
rect 2094 4162 2124 4171
rect 2106 4160 2124 4162
rect 2161 4144 2167 4228
rect 2273 4232 2279 4246
rect 2321 4238 2327 4256
rect 2235 4226 2279 4232
rect 2287 4232 2327 4238
rect 2206 4187 2233 4194
rect 2180 4176 2186 4181
rect 2180 4168 2214 4176
rect 2219 4160 2226 4168
rect 2287 4160 2293 4232
rect 2347 4224 2361 4232
rect 2353 4173 2367 4187
rect 2375 4173 2383 4236
rect 2397 4230 2405 4276
rect 2397 4224 2423 4230
rect 2420 4218 2423 4224
rect 2219 4154 2293 4160
rect 2367 4159 2383 4173
rect 2219 4148 2226 4154
rect 2287 4152 2293 4154
rect 2251 4136 2272 4143
rect 2375 4144 2383 4159
rect 2420 4162 2427 4218
rect 2441 4201 2449 4236
rect 2447 4187 2449 4201
rect 2496 4193 2504 4276
rect 2667 4262 2679 4296
rect 2721 4270 2733 4276
rect 2775 4270 2783 4276
rect 2725 4258 2747 4270
rect 2775 4256 2793 4270
rect 2673 4238 2679 4256
rect 2697 4246 2727 4252
rect 2775 4250 2783 4256
rect 2563 4229 2580 4236
rect 2420 4156 2423 4162
rect 2200 4124 2207 4130
rect 2265 4124 2272 4136
rect 2322 4130 2333 4138
rect 2322 4124 2329 4130
rect 2200 4118 2213 4124
rect 2401 4150 2423 4156
rect 2401 4124 2409 4150
rect 2441 4144 2449 4187
rect 2573 4181 2580 4229
rect 2496 4124 2504 4179
rect 2617 4173 2625 4236
rect 2639 4224 2653 4232
rect 2673 4232 2713 4238
rect 2633 4173 2647 4187
rect 2573 4124 2580 4167
rect 2617 4159 2633 4173
rect 2707 4160 2713 4232
rect 2721 4232 2727 4246
rect 2745 4242 2783 4250
rect 2721 4226 2765 4232
rect 2777 4228 2839 4236
rect 2767 4187 2794 4194
rect 2814 4176 2820 4181
rect 2786 4168 2820 4176
rect 2774 4160 2781 4168
rect 2617 4144 2625 4159
rect 2707 4154 2781 4160
rect 2707 4152 2713 4154
rect 1897 4098 1909 4104
rect 1958 4098 1970 4104
rect 2058 4098 2070 4104
rect 2181 4098 2193 4104
rect 2243 4098 2255 4104
rect 2291 4098 2303 4104
rect 2349 4098 2361 4104
rect 2419 4098 2431 4104
rect 2511 4098 2523 4104
rect 2774 4148 2781 4154
rect 2667 4130 2678 4138
rect 2671 4124 2678 4130
rect 2728 4136 2749 4143
rect 2833 4144 2839 4228
rect 2876 4193 2884 4276
rect 3002 4316 3014 4322
rect 3052 4316 3064 4322
rect 3097 4316 3109 4322
rect 3137 4316 3149 4322
rect 3191 4316 3203 4322
rect 3231 4316 3243 4322
rect 3271 4316 3283 4322
rect 3311 4316 3323 4322
rect 3337 4316 3349 4322
rect 3441 4316 3453 4322
rect 3507 4316 3519 4322
rect 3553 4316 3565 4322
rect 3611 4316 3623 4322
rect 3671 4316 3683 4322
rect 3711 4316 3723 4322
rect 2943 4229 2960 4236
rect 2953 4181 2960 4229
rect 3033 4201 3041 4236
rect 3117 4221 3125 4276
rect 3215 4221 3223 4276
rect 3295 4221 3303 4276
rect 3360 4229 3377 4236
rect 3477 4270 3485 4276
rect 3527 4270 3539 4276
rect 3467 4256 3485 4270
rect 3513 4258 3535 4270
rect 3581 4262 3593 4296
rect 3477 4250 3485 4256
rect 3477 4242 3515 4250
rect 3533 4246 3563 4252
rect 2728 4124 2735 4136
rect 2793 4124 2800 4130
rect 2787 4118 2800 4124
rect 2876 4124 2884 4179
rect 2953 4124 2960 4167
rect 3039 4165 3047 4187
rect 3040 4158 3065 4165
rect 2997 4144 3049 4147
rect 3009 4138 3037 4144
rect 3057 4144 3065 4158
rect 3117 4158 3125 4207
rect 3215 4158 3223 4207
rect 3295 4158 3303 4207
rect 3360 4181 3367 4229
rect 3421 4228 3483 4236
rect 3117 4152 3141 4158
rect 3129 4144 3141 4152
rect 3199 4152 3223 4158
rect 3279 4152 3303 4158
rect 3199 4144 3211 4152
rect 3279 4144 3291 4152
rect 3360 4124 3367 4167
rect 3421 4144 3427 4228
rect 3533 4232 3539 4246
rect 3581 4238 3587 4256
rect 3495 4226 3539 4232
rect 3547 4232 3587 4238
rect 3466 4187 3493 4194
rect 3440 4176 3446 4181
rect 3440 4168 3474 4176
rect 3479 4160 3486 4168
rect 3547 4160 3553 4232
rect 3737 4316 3749 4322
rect 3837 4316 3849 4322
rect 3895 4316 3907 4322
rect 3941 4316 3953 4322
rect 4007 4316 4019 4322
rect 4057 4316 4069 4322
rect 4191 4316 4203 4322
rect 4259 4316 4271 4322
rect 4371 4316 4383 4322
rect 4451 4316 4463 4322
rect 4517 4316 4529 4322
rect 4575 4316 4587 4322
rect 4621 4316 4633 4322
rect 4687 4316 4699 4322
rect 3607 4224 3621 4232
rect 3613 4173 3627 4187
rect 3635 4173 3643 4236
rect 3695 4221 3703 4276
rect 3760 4229 3777 4236
rect 3867 4262 3879 4296
rect 3921 4270 3933 4276
rect 3975 4270 3983 4276
rect 3925 4258 3947 4270
rect 3975 4256 3993 4270
rect 3873 4238 3879 4256
rect 3897 4246 3927 4252
rect 3975 4250 3983 4256
rect 3479 4154 3553 4160
rect 3627 4159 3643 4173
rect 3479 4148 3486 4154
rect 3547 4152 3553 4154
rect 2551 4098 2563 4104
rect 2591 4098 2603 4104
rect 2639 4098 2651 4104
rect 2697 4098 2709 4104
rect 2745 4098 2757 4104
rect 2807 4098 2819 4104
rect 2857 4098 2869 4104
rect 2931 4098 2943 4104
rect 2971 4098 2983 4104
rect 3017 4098 3029 4104
rect 3099 4098 3111 4104
rect 3229 4098 3241 4104
rect 3309 4098 3321 4104
rect 3511 4136 3532 4143
rect 3635 4144 3643 4159
rect 3695 4158 3703 4207
rect 3760 4181 3767 4229
rect 3460 4124 3467 4130
rect 3525 4124 3532 4136
rect 3582 4130 3593 4138
rect 3582 4124 3589 4130
rect 3460 4118 3473 4124
rect 3679 4152 3703 4158
rect 3679 4144 3691 4152
rect 3760 4124 3767 4167
rect 3817 4173 3825 4236
rect 3839 4224 3853 4232
rect 3873 4232 3913 4238
rect 3833 4173 3847 4187
rect 3817 4159 3833 4173
rect 3907 4160 3913 4232
rect 3921 4232 3927 4246
rect 3945 4242 3983 4250
rect 4211 4242 4223 4244
rect 4183 4236 4223 4242
rect 3921 4226 3965 4232
rect 3977 4228 4039 4236
rect 3967 4187 3994 4194
rect 4014 4176 4020 4181
rect 3986 4168 4020 4176
rect 3974 4160 3981 4168
rect 3817 4144 3825 4159
rect 3907 4154 3981 4160
rect 3907 4152 3913 4154
rect 3337 4098 3349 4104
rect 3377 4098 3389 4104
rect 3441 4098 3453 4104
rect 3503 4098 3515 4104
rect 3551 4098 3563 4104
rect 3609 4098 3621 4104
rect 3709 4098 3721 4104
rect 3974 4148 3981 4154
rect 3867 4130 3878 4138
rect 3871 4124 3878 4130
rect 3928 4136 3949 4143
rect 4033 4144 4039 4228
rect 4080 4229 4097 4236
rect 4080 4181 4087 4229
rect 4154 4201 4162 4236
rect 4237 4230 4245 4276
rect 4471 4242 4483 4244
rect 4443 4236 4483 4242
rect 4547 4262 4559 4296
rect 4601 4270 4613 4276
rect 4655 4270 4663 4276
rect 4605 4258 4627 4270
rect 4655 4256 4673 4270
rect 4553 4238 4559 4256
rect 4577 4246 4607 4252
rect 4655 4250 4663 4256
rect 4237 4224 4263 4230
rect 4260 4218 4263 4224
rect 3928 4124 3935 4136
rect 3993 4124 4000 4130
rect 3987 4118 4000 4124
rect 4080 4124 4087 4167
rect 4154 4144 4162 4187
rect 4260 4162 4267 4218
rect 4281 4201 4289 4236
rect 4343 4229 4360 4236
rect 4287 4187 4289 4201
rect 4260 4156 4263 4162
rect 4241 4150 4263 4156
rect 4154 4133 4180 4144
rect 3737 4098 3749 4104
rect 3777 4098 3789 4104
rect 3839 4098 3851 4104
rect 3897 4098 3909 4104
rect 3945 4098 3957 4104
rect 4007 4098 4019 4104
rect 4057 4098 4069 4104
rect 4097 4098 4109 4104
rect 4241 4124 4249 4150
rect 4281 4144 4289 4187
rect 4353 4181 4360 4229
rect 4414 4201 4422 4236
rect 4353 4124 4360 4167
rect 4414 4144 4422 4187
rect 4497 4173 4505 4236
rect 4519 4224 4533 4232
rect 4553 4232 4593 4238
rect 4513 4173 4527 4187
rect 4497 4159 4513 4173
rect 4587 4160 4593 4232
rect 4601 4232 4607 4246
rect 4625 4242 4663 4250
rect 4601 4226 4645 4232
rect 4657 4228 4719 4236
rect 4647 4187 4674 4194
rect 4694 4176 4700 4181
rect 4666 4168 4700 4176
rect 4654 4160 4661 4168
rect 4497 4144 4505 4159
rect 4587 4154 4661 4160
rect 4587 4152 4593 4154
rect 4414 4133 4440 4144
rect 4158 4098 4170 4104
rect 4208 4098 4220 4104
rect 4259 4098 4271 4104
rect 4331 4098 4343 4104
rect 4371 4098 4383 4104
rect 4654 4148 4661 4154
rect 4547 4130 4558 4138
rect 4551 4124 4558 4130
rect 4608 4136 4629 4143
rect 4713 4144 4719 4228
rect 4608 4124 4615 4136
rect 4673 4124 4680 4130
rect 4667 4118 4680 4124
rect 4418 4098 4430 4104
rect 4468 4098 4480 4104
rect 4519 4098 4531 4104
rect 4577 4098 4589 4104
rect 4625 4098 4637 4104
rect 4687 4098 4699 4104
rect 4782 4098 4842 4562
rect 4 4096 4842 4098
rect 4776 4084 4842 4096
rect 4 4082 4842 4084
rect 69 4076 81 4082
rect 99 4076 111 4082
rect 229 4076 241 4082
rect 311 4076 323 4082
rect 360 4076 372 4082
rect 410 4076 422 4082
rect 39 4028 51 4036
rect 129 4028 141 4036
rect 39 4022 63 4028
rect 55 3973 63 4022
rect 117 4022 141 4028
rect 199 4028 211 4036
rect 199 4022 223 4028
rect 117 3973 125 4022
rect 215 3973 223 4022
rect 275 4022 283 4036
rect 303 4036 331 4042
rect 471 4076 483 4082
rect 511 4076 523 4082
rect 539 4076 551 4082
rect 637 4076 649 4082
rect 790 4076 802 4082
rect 400 4036 426 4047
rect 291 4033 343 4036
rect 275 4015 300 4022
rect 293 3993 301 4015
rect 418 3993 426 4036
rect 493 4013 500 4056
rect 569 4028 581 4036
rect 629 4036 657 4042
rect 617 4033 669 4036
rect 557 4022 581 4028
rect 677 4022 685 4036
rect 55 3904 63 3959
rect 117 3904 125 3959
rect 215 3904 223 3959
rect 299 3944 307 3979
rect 418 3944 426 3979
rect 493 3951 500 3999
rect 557 3973 565 4022
rect 660 4015 685 4022
rect 736 4018 754 4020
rect 659 3993 667 4015
rect 736 4009 766 4018
rect 818 4076 830 4082
rect 971 4076 983 4082
rect 1037 4076 1049 4082
rect 1151 4076 1163 4082
rect 1250 4076 1262 4082
rect 935 4022 943 4036
rect 963 4036 991 4042
rect 951 4033 1003 4036
rect 1029 4036 1057 4042
rect 1017 4033 1069 4036
rect 1077 4022 1085 4036
rect 866 4018 884 4020
rect 854 4009 884 4018
rect 935 4015 960 4022
rect 1060 4015 1085 4022
rect 736 3981 744 4009
rect 876 3981 884 4009
rect 953 3993 961 4015
rect 483 3944 500 3951
rect 31 3858 43 3864
rect 71 3858 83 3864
rect 97 3858 109 3864
rect 137 3858 149 3864
rect 191 3858 203 3864
rect 231 3858 243 3864
rect 357 3938 397 3944
rect 357 3936 369 3938
rect 557 3904 565 3959
rect 653 3944 661 3979
rect 276 3858 288 3864
rect 326 3858 338 3864
rect 377 3858 389 3864
rect 511 3858 523 3864
rect 537 3858 549 3864
rect 577 3858 589 3864
rect 735 3912 742 3967
rect 1059 3993 1067 4015
rect 1136 4001 1144 4056
rect 1196 4018 1214 4020
rect 1196 4009 1226 4018
rect 1277 4076 1289 4082
rect 1338 4076 1350 4082
rect 1438 4076 1450 4082
rect 1539 4076 1551 4082
rect 1631 4076 1643 4082
rect 1671 4076 1683 4082
rect 1741 4076 1753 4082
rect 1851 4076 1863 4082
rect 1897 4076 1909 4082
rect 1937 4076 1949 4082
rect 2011 4076 2023 4082
rect 2057 4076 2069 4082
rect 2137 4076 2149 4082
rect 2199 4076 2211 4082
rect 2278 4076 2290 4082
rect 2399 4076 2411 4082
rect 2457 4076 2469 4082
rect 2497 4076 2509 4082
rect 2537 4076 2549 4082
rect 2577 4076 2589 4082
rect 2617 4076 2629 4082
rect 2681 4076 2693 4082
rect 2743 4076 2755 4082
rect 2791 4076 2803 4082
rect 2849 4076 2861 4082
rect 2897 4076 2909 4082
rect 2977 4076 2989 4082
rect 3057 4076 3069 4082
rect 3097 4076 3109 4082
rect 878 3912 885 3967
rect 959 3944 967 3979
rect 1053 3944 1061 3979
rect 735 3906 782 3912
rect 735 3904 743 3906
rect 771 3904 782 3906
rect 838 3906 885 3912
rect 838 3904 849 3906
rect 622 3858 634 3864
rect 672 3858 684 3864
rect 751 3858 763 3864
rect 791 3858 803 3864
rect 877 3904 885 3906
rect 817 3858 829 3864
rect 857 3858 869 3864
rect 936 3858 948 3864
rect 986 3858 998 3864
rect 1136 3904 1144 3987
rect 1196 3981 1204 4009
rect 1296 4001 1304 4056
rect 1386 4018 1404 4020
rect 1374 4009 1404 4018
rect 1569 4028 1581 4036
rect 1557 4022 1581 4028
rect 1486 4018 1504 4020
rect 1474 4009 1504 4018
rect 1195 3912 1202 3967
rect 1195 3906 1242 3912
rect 1195 3904 1203 3906
rect 1231 3904 1242 3906
rect 1296 3904 1304 3987
rect 1396 3981 1404 4009
rect 1496 3981 1504 4009
rect 1398 3912 1405 3967
rect 1557 3973 1565 4022
rect 1653 4013 1660 4056
rect 1711 4036 1721 4046
rect 1498 3912 1505 3967
rect 1358 3906 1405 3912
rect 1358 3904 1369 3906
rect 1022 3858 1034 3864
rect 1072 3858 1084 3864
rect 1151 3858 1163 3864
rect 1211 3858 1223 3864
rect 1251 3858 1263 3864
rect 1397 3904 1405 3906
rect 1458 3906 1505 3912
rect 1458 3904 1469 3906
rect 1497 3904 1505 3906
rect 1557 3904 1565 3959
rect 1653 3951 1660 3999
rect 1711 3993 1719 4036
rect 1771 4026 1783 4036
rect 1745 4018 1783 4026
rect 1815 4022 1823 4036
rect 1843 4036 1871 4042
rect 1831 4033 1883 4036
rect 1711 3979 1713 3993
rect 1643 3944 1660 3951
rect 1711 3944 1719 3979
rect 1754 3904 1762 4018
rect 1815 4015 1840 4022
rect 1833 3993 1841 4015
rect 1920 4013 1927 4056
rect 1996 4001 2004 4056
rect 2049 4036 2077 4042
rect 2037 4033 2089 4036
rect 2097 4022 2105 4036
rect 2080 4015 2105 4022
rect 1839 3944 1847 3979
rect 1920 3951 1927 3999
rect 1920 3944 1937 3951
rect 1277 3858 1289 3864
rect 1337 3858 1349 3864
rect 1377 3858 1389 3864
rect 1437 3858 1449 3864
rect 1477 3858 1489 3864
rect 1537 3858 1549 3864
rect 1577 3858 1589 3864
rect 1671 3858 1683 3864
rect 1727 3858 1739 3864
rect 1771 3858 1783 3864
rect 1816 3858 1828 3864
rect 1866 3858 1878 3864
rect 1996 3904 2004 3987
rect 2079 3993 2087 4015
rect 2156 4001 2164 4056
rect 2229 4028 2241 4036
rect 2217 4022 2241 4028
rect 2073 3944 2081 3979
rect 1897 3858 1909 3864
rect 2011 3858 2023 3864
rect 2156 3904 2164 3987
rect 2217 3973 2225 4022
rect 2381 4030 2389 4056
rect 2700 4056 2713 4062
rect 2700 4050 2707 4056
rect 2765 4044 2772 4056
rect 2381 4024 2403 4030
rect 2326 4018 2344 4020
rect 2314 4009 2344 4018
rect 2336 3981 2344 4009
rect 2400 4018 2403 4024
rect 2217 3904 2225 3959
rect 2338 3912 2345 3967
rect 2400 3962 2407 4018
rect 2421 3993 2429 4036
rect 2476 4030 2488 4036
rect 2517 4030 2529 4036
rect 2556 4030 2568 4036
rect 2596 4030 2608 4036
rect 2476 4022 2503 4030
rect 2517 4022 2542 4030
rect 2556 4022 2582 4030
rect 2596 4029 2614 4030
rect 2596 4022 2615 4029
rect 2495 4016 2503 4022
rect 2534 4016 2542 4022
rect 2574 4016 2582 4022
rect 2495 4004 2510 4016
rect 2534 4004 2550 4016
rect 2574 4004 2590 4016
rect 2427 3979 2429 3993
rect 2400 3956 2403 3962
rect 2298 3906 2345 3912
rect 2298 3904 2309 3906
rect 2042 3858 2054 3864
rect 2092 3858 2104 3864
rect 2137 3858 2149 3864
rect 2197 3858 2209 3864
rect 2237 3858 2249 3864
rect 2337 3904 2345 3906
rect 2377 3950 2403 3956
rect 2377 3904 2385 3950
rect 2421 3944 2429 3979
rect 2495 3958 2503 4004
rect 2534 3958 2542 4004
rect 2574 3958 2582 4004
rect 2608 4001 2615 4022
rect 2608 3987 2613 4001
rect 2608 3958 2615 3987
rect 2477 3950 2503 3958
rect 2517 3950 2542 3958
rect 2557 3950 2582 3958
rect 2597 3950 2615 3958
rect 2661 3952 2667 4036
rect 2751 4037 2772 4044
rect 2822 4050 2829 4056
rect 2822 4042 2833 4050
rect 2719 4026 2726 4032
rect 2787 4026 2793 4028
rect 2719 4020 2793 4026
rect 2875 4021 2883 4036
rect 2719 4012 2726 4020
rect 2680 4004 2714 4012
rect 2680 3999 2686 4004
rect 2706 3986 2733 3993
rect 2477 3944 2489 3950
rect 2517 3944 2529 3950
rect 2557 3944 2569 3950
rect 2597 3944 2609 3950
rect 2661 3944 2723 3952
rect 2735 3948 2779 3954
rect 2717 3930 2755 3938
rect 2773 3934 2779 3948
rect 2787 3948 2793 4020
rect 2867 4007 2883 4021
rect 2853 3993 2867 4007
rect 2787 3942 2827 3948
rect 2847 3948 2861 3956
rect 2875 3944 2883 4007
rect 2916 4001 2924 4056
rect 2969 4036 2997 4042
rect 2957 4033 3009 4036
rect 3139 4076 3151 4082
rect 3238 4076 3250 4082
rect 3288 4076 3300 4082
rect 3347 4076 3359 4082
rect 3431 4076 3443 4082
rect 3471 4076 3483 4082
rect 3531 4076 3543 4082
rect 3579 4076 3591 4082
rect 3637 4076 3649 4082
rect 3685 4076 3697 4082
rect 3747 4076 3759 4082
rect 3818 4076 3830 4082
rect 3868 4076 3880 4082
rect 3017 4022 3025 4036
rect 3000 4015 3025 4022
rect 2717 3924 2725 3930
rect 2773 3928 2803 3934
rect 2821 3924 2827 3942
rect 2707 3910 2725 3924
rect 2753 3910 2775 3922
rect 2717 3904 2725 3910
rect 2767 3904 2779 3910
rect 2821 3884 2833 3918
rect 2916 3904 2924 3987
rect 2999 3993 3007 4015
rect 3080 4013 3087 4056
rect 3169 4028 3181 4036
rect 2993 3944 3001 3979
rect 3080 3951 3087 3999
rect 3157 4022 3181 4028
rect 3234 4036 3260 4047
rect 3379 4036 3389 4046
rect 3157 3973 3165 4022
rect 3234 3993 3242 4036
rect 3317 4026 3329 4036
rect 3317 4018 3355 4026
rect 3080 3944 3097 3951
rect 2277 3858 2289 3864
rect 2317 3858 2329 3864
rect 2399 3858 2411 3864
rect 2457 3858 2469 3864
rect 2497 3858 2509 3864
rect 2537 3858 2549 3864
rect 2577 3858 2589 3864
rect 2617 3858 2629 3864
rect 2681 3858 2693 3864
rect 2747 3858 2759 3864
rect 2793 3858 2805 3864
rect 2851 3858 2863 3864
rect 2897 3858 2909 3864
rect 2962 3858 2974 3864
rect 3012 3858 3024 3864
rect 3157 3904 3165 3959
rect 3234 3944 3242 3979
rect 3263 3938 3303 3944
rect 3291 3936 3303 3938
rect 3338 3904 3346 4018
rect 3381 3993 3389 4036
rect 3453 4013 3460 4056
rect 3516 4001 3524 4056
rect 3727 4056 3740 4062
rect 3611 4050 3618 4056
rect 3607 4042 3618 4050
rect 3668 4044 3675 4056
rect 3733 4050 3740 4056
rect 3557 4021 3565 4036
rect 3668 4037 3689 4044
rect 3647 4026 3653 4028
rect 3714 4026 3721 4032
rect 3387 3979 3389 3993
rect 3381 3944 3389 3979
rect 3453 3951 3460 3999
rect 3557 4007 3573 4021
rect 3647 4020 3721 4026
rect 3443 3944 3460 3951
rect 3516 3904 3524 3987
rect 3557 3944 3565 4007
rect 3573 3993 3587 4007
rect 3579 3948 3593 3956
rect 3647 3948 3653 4020
rect 3714 4012 3721 4020
rect 3726 4004 3760 4012
rect 3754 3999 3760 4004
rect 3707 3986 3734 3993
rect 3613 3942 3653 3948
rect 3661 3948 3705 3954
rect 3613 3924 3619 3942
rect 3661 3934 3667 3948
rect 3773 3952 3779 4036
rect 3814 4036 3840 4047
rect 3897 4076 3909 4082
rect 3937 4076 3949 4082
rect 3991 4076 4003 4082
rect 4031 4076 4043 4082
rect 4087 4076 4099 4082
rect 4177 4076 4189 4082
rect 4311 4076 4323 4082
rect 4391 4076 4403 4082
rect 4439 4076 4451 4082
rect 4497 4076 4509 4082
rect 4545 4076 4557 4082
rect 4607 4076 4619 4082
rect 4657 4076 4669 4082
rect 3814 3993 3822 4036
rect 3920 4013 3927 4056
rect 3717 3944 3779 3952
rect 3814 3944 3822 3979
rect 3920 3951 3927 3999
rect 4013 4013 4020 4056
rect 4119 4036 4129 4046
rect 4057 4026 4069 4036
rect 4057 4018 4095 4026
rect 4013 3951 4020 3999
rect 3920 3944 3937 3951
rect 3637 3928 3667 3934
rect 3685 3930 3723 3938
rect 3715 3924 3723 3930
rect 3607 3884 3619 3918
rect 3665 3910 3687 3922
rect 3715 3910 3733 3924
rect 3661 3904 3673 3910
rect 3715 3904 3723 3910
rect 3843 3938 3883 3944
rect 3871 3936 3883 3938
rect 4003 3944 4020 3951
rect 4078 3904 4086 4018
rect 4121 3993 4129 4036
rect 4169 4036 4197 4042
rect 4157 4033 4209 4036
rect 4217 4022 4225 4036
rect 4200 4015 4225 4022
rect 4275 4022 4283 4036
rect 4303 4036 4331 4042
rect 4291 4033 4343 4036
rect 4275 4015 4300 4022
rect 4127 3979 4129 3993
rect 4199 3993 4207 4015
rect 4293 3993 4301 4015
rect 4347 4017 4363 4023
rect 4121 3944 4129 3979
rect 4193 3944 4201 3979
rect 4299 3944 4307 3979
rect 4357 3967 4363 4017
rect 4376 4001 4384 4056
rect 4587 4056 4600 4062
rect 4471 4050 4478 4056
rect 4467 4042 4478 4050
rect 4528 4044 4535 4056
rect 4593 4050 4600 4056
rect 4417 4021 4425 4036
rect 4528 4037 4549 4044
rect 4507 4026 4513 4028
rect 4574 4026 4581 4032
rect 4417 4007 4433 4021
rect 4507 4020 4581 4026
rect 3057 3858 3069 3864
rect 3137 3858 3149 3864
rect 3177 3858 3189 3864
rect 3271 3858 3283 3864
rect 3317 3858 3329 3864
rect 3361 3858 3373 3864
rect 3471 3858 3483 3864
rect 3531 3858 3543 3864
rect 3577 3858 3589 3864
rect 3635 3858 3647 3864
rect 3681 3858 3693 3864
rect 3747 3858 3759 3864
rect 3851 3858 3863 3864
rect 3897 3858 3909 3864
rect 4031 3858 4043 3864
rect 4057 3858 4069 3864
rect 4101 3858 4113 3864
rect 4162 3858 4174 3864
rect 4212 3858 4224 3864
rect 4376 3904 4384 3987
rect 4417 3944 4425 4007
rect 4433 3993 4447 4007
rect 4439 3948 4453 3956
rect 4507 3948 4513 4020
rect 4574 4012 4581 4020
rect 4586 4004 4620 4012
rect 4614 3999 4620 4004
rect 4567 3986 4594 3993
rect 4473 3942 4513 3948
rect 4521 3948 4565 3954
rect 4473 3924 4479 3942
rect 4521 3934 4527 3948
rect 4633 3952 4639 4036
rect 4676 4001 4684 4056
rect 4577 3944 4639 3952
rect 4497 3928 4527 3934
rect 4545 3930 4583 3938
rect 4575 3924 4583 3930
rect 4467 3884 4479 3918
rect 4525 3910 4547 3922
rect 4575 3910 4593 3924
rect 4521 3904 4533 3910
rect 4575 3904 4583 3910
rect 4676 3904 4684 3987
rect 4276 3858 4288 3864
rect 4326 3858 4338 3864
rect 4391 3858 4403 3864
rect 4437 3858 4449 3864
rect 4495 3858 4507 3864
rect 4541 3858 4553 3864
rect 4607 3858 4619 3864
rect 4657 3858 4669 3864
rect -62 3856 4776 3858
rect -62 3844 4 3856
rect -62 3842 4776 3844
rect -62 3378 -2 3842
rect 71 3836 83 3842
rect 102 3836 114 3842
rect 152 3836 164 3842
rect 231 3836 243 3842
rect 311 3836 323 3842
rect 387 3836 399 3842
rect 431 3836 443 3842
rect 43 3749 60 3756
rect 53 3701 60 3749
rect 133 3721 141 3756
rect 216 3713 224 3796
rect 331 3762 343 3764
rect 303 3756 343 3762
rect 471 3836 483 3842
rect 511 3836 523 3842
rect 551 3836 563 3842
rect 591 3836 603 3842
rect 617 3836 629 3842
rect 682 3836 694 3842
rect 732 3836 744 3842
rect 274 3721 282 3756
rect 371 3721 379 3756
rect 53 3644 60 3687
rect 139 3685 147 3707
rect 140 3678 165 3685
rect 97 3664 149 3667
rect 109 3658 137 3664
rect 157 3664 165 3678
rect 216 3644 224 3699
rect 274 3664 282 3707
rect 371 3707 373 3721
rect 371 3664 379 3707
rect 414 3682 422 3796
rect 495 3741 503 3796
rect 537 3757 553 3763
rect 405 3674 443 3682
rect 495 3678 503 3727
rect 537 3687 543 3757
rect 575 3741 583 3796
rect 431 3664 443 3674
rect 274 3653 300 3664
rect 31 3618 43 3624
rect 71 3618 83 3624
rect 117 3618 129 3624
rect 231 3618 243 3624
rect 371 3654 381 3664
rect 479 3672 503 3678
rect 575 3678 583 3727
rect 636 3713 644 3796
rect 777 3836 789 3842
rect 817 3836 829 3842
rect 891 3836 903 3842
rect 931 3836 943 3842
rect 977 3836 989 3842
rect 1057 3836 1069 3842
rect 1097 3836 1109 3842
rect 1177 3836 1189 3842
rect 1257 3836 1269 3842
rect 1351 3836 1363 3842
rect 1391 3836 1403 3842
rect 1451 3836 1463 3842
rect 713 3721 721 3756
rect 559 3672 583 3678
rect 479 3664 491 3672
rect 559 3664 571 3672
rect 636 3644 644 3699
rect 719 3685 727 3707
rect 757 3703 763 3753
rect 797 3741 805 3796
rect 875 3794 883 3796
rect 911 3794 922 3796
rect 875 3788 922 3794
rect 875 3733 882 3788
rect 957 3762 969 3764
rect 957 3756 997 3762
rect 1078 3794 1089 3796
rect 1117 3794 1125 3796
rect 1078 3788 1125 3794
rect 747 3697 763 3703
rect 720 3678 745 3685
rect 677 3664 729 3667
rect 278 3618 290 3624
rect 328 3618 340 3624
rect 401 3618 413 3624
rect 509 3618 521 3624
rect 589 3618 601 3624
rect 689 3658 717 3664
rect 737 3664 745 3678
rect 797 3678 805 3727
rect 1018 3721 1026 3756
rect 1118 3733 1125 3788
rect 1157 3762 1169 3764
rect 1157 3756 1197 3762
rect 876 3691 884 3719
rect 876 3682 906 3691
rect 1218 3721 1226 3756
rect 876 3680 894 3682
rect 797 3672 821 3678
rect 809 3664 821 3672
rect 1018 3664 1026 3707
rect 1116 3691 1124 3719
rect 617 3618 629 3624
rect 697 3618 709 3624
rect 779 3618 791 3624
rect 930 3618 942 3624
rect 1000 3653 1026 3664
rect 960 3618 972 3624
rect 1010 3618 1022 3624
rect 1094 3682 1124 3691
rect 1276 3713 1284 3796
rect 1335 3794 1343 3796
rect 1496 3836 1508 3842
rect 1546 3836 1558 3842
rect 1611 3836 1623 3842
rect 1657 3836 1669 3842
rect 1737 3836 1749 3842
rect 1871 3836 1883 3842
rect 1931 3836 1943 3842
rect 1971 3836 1983 3842
rect 2027 3836 2039 3842
rect 2119 3836 2131 3842
rect 2191 3836 2203 3842
rect 2231 3836 2243 3842
rect 2271 3836 2283 3842
rect 2311 3836 2323 3842
rect 2351 3836 2363 3842
rect 2401 3836 2413 3842
rect 2467 3836 2479 3842
rect 2513 3836 2525 3842
rect 2571 3836 2583 3842
rect 2636 3836 2648 3842
rect 2686 3836 2698 3842
rect 2751 3836 2763 3842
rect 2831 3836 2843 3842
rect 2911 3836 2923 3842
rect 2991 3836 3003 3842
rect 1371 3794 1382 3796
rect 1335 3788 1382 3794
rect 1335 3733 1342 3788
rect 1106 3680 1124 3682
rect 1218 3664 1226 3707
rect 1200 3653 1226 3664
rect 1276 3644 1284 3699
rect 1336 3691 1344 3719
rect 1436 3713 1444 3796
rect 1519 3721 1527 3756
rect 1336 3682 1366 3691
rect 1336 3680 1354 3682
rect 1058 3618 1070 3624
rect 1160 3618 1172 3624
rect 1210 3618 1222 3624
rect 1436 3644 1444 3699
rect 1513 3685 1521 3707
rect 1596 3713 1604 3796
rect 1637 3762 1649 3764
rect 1637 3756 1677 3762
rect 1891 3762 1903 3764
rect 1863 3756 1903 3762
rect 1698 3721 1706 3756
rect 1760 3749 1777 3756
rect 1495 3678 1520 3685
rect 1495 3664 1503 3678
rect 1511 3664 1563 3667
rect 1523 3658 1551 3664
rect 1596 3644 1604 3699
rect 1698 3664 1706 3707
rect 1760 3701 1767 3749
rect 1834 3721 1842 3756
rect 1955 3741 1963 3796
rect 2059 3757 2063 3766
rect 1997 3748 2005 3756
rect 1997 3740 2033 3748
rect 1257 3618 1269 3624
rect 1390 3618 1402 3624
rect 1451 3618 1463 3624
rect 1531 3618 1543 3624
rect 1611 3618 1623 3624
rect 1680 3653 1706 3664
rect 1760 3644 1767 3687
rect 1834 3664 1842 3707
rect 1955 3678 1963 3727
rect 2038 3684 2044 3739
rect 2054 3713 2063 3757
rect 2097 3750 2105 3796
rect 2437 3790 2445 3796
rect 2487 3790 2499 3796
rect 2427 3776 2445 3790
rect 2473 3778 2495 3790
rect 2541 3782 2553 3816
rect 2437 3770 2445 3776
rect 2437 3762 2475 3770
rect 2493 3766 2523 3772
rect 2097 3744 2123 3750
rect 2120 3738 2123 3744
rect 1939 3672 1963 3678
rect 2023 3672 2033 3678
rect 1939 3664 1951 3672
rect 1834 3653 1860 3664
rect 1640 3618 1652 3624
rect 1690 3618 1702 3624
rect 1737 3618 1749 3624
rect 1777 3618 1789 3624
rect 2023 3644 2029 3672
rect 2060 3664 2067 3699
rect 2120 3682 2127 3738
rect 2141 3721 2149 3756
rect 2211 3750 2223 3756
rect 2251 3750 2263 3756
rect 2291 3750 2303 3756
rect 2331 3750 2343 3756
rect 2147 3707 2149 3721
rect 2205 3742 2223 3750
rect 2238 3742 2263 3750
rect 2278 3742 2303 3750
rect 2317 3742 2343 3750
rect 2381 3748 2443 3756
rect 2205 3713 2212 3742
rect 2120 3676 2123 3682
rect 2101 3670 2123 3676
rect 1838 3618 1850 3624
rect 1888 3618 1900 3624
rect 1969 3618 1981 3624
rect 2101 3644 2109 3670
rect 2141 3664 2149 3707
rect 2207 3699 2212 3713
rect 2205 3678 2212 3699
rect 2238 3696 2246 3742
rect 2278 3696 2286 3742
rect 2317 3696 2325 3742
rect 2230 3684 2246 3696
rect 2270 3684 2286 3696
rect 2310 3684 2325 3696
rect 2238 3678 2246 3684
rect 2278 3678 2286 3684
rect 2317 3678 2325 3684
rect 2205 3671 2224 3678
rect 2206 3670 2224 3671
rect 2238 3670 2264 3678
rect 2278 3670 2303 3678
rect 2317 3670 2344 3678
rect 2212 3664 2224 3670
rect 2252 3664 2264 3670
rect 2291 3664 2303 3670
rect 2332 3664 2344 3670
rect 2381 3664 2387 3748
rect 2493 3752 2499 3766
rect 2541 3758 2547 3776
rect 2455 3746 2499 3752
rect 2507 3752 2547 3758
rect 2426 3707 2453 3714
rect 2400 3696 2406 3701
rect 2400 3688 2434 3696
rect 2439 3680 2446 3688
rect 2507 3680 2513 3752
rect 2567 3744 2581 3752
rect 2573 3693 2587 3707
rect 2595 3693 2603 3756
rect 2659 3721 2667 3756
rect 2439 3674 2513 3680
rect 2587 3679 2603 3693
rect 2653 3685 2661 3707
rect 2736 3713 2744 3796
rect 3017 3836 3029 3842
rect 3111 3836 3123 3842
rect 3142 3836 3154 3842
rect 3192 3836 3204 3842
rect 3291 3836 3303 3842
rect 3357 3836 3369 3842
rect 3437 3836 3449 3842
rect 3497 3836 3509 3842
rect 3541 3836 3553 3842
rect 3602 3836 3614 3842
rect 3652 3836 3664 3842
rect 2803 3749 2820 3756
rect 2883 3749 2900 3756
rect 2963 3749 2980 3756
rect 2813 3701 2820 3749
rect 2893 3701 2900 3749
rect 2973 3701 2980 3749
rect 3036 3713 3044 3796
rect 3096 3713 3104 3796
rect 3311 3762 3323 3764
rect 3283 3756 3323 3762
rect 3337 3762 3349 3764
rect 3337 3756 3377 3762
rect 3173 3721 3181 3756
rect 3254 3721 3262 3756
rect 3398 3721 3406 3756
rect 2439 3668 2446 3674
rect 2507 3672 2513 3674
rect 2471 3656 2492 3663
rect 2595 3664 2603 3679
rect 2635 3678 2660 3685
rect 2635 3664 2643 3678
rect 2420 3644 2427 3650
rect 2485 3644 2492 3656
rect 2542 3650 2553 3658
rect 2542 3644 2549 3650
rect 2420 3638 2433 3644
rect 2651 3664 2703 3667
rect 2663 3658 2691 3664
rect 2736 3644 2744 3699
rect 2813 3644 2820 3687
rect 2893 3644 2900 3687
rect 2973 3644 2980 3687
rect 3036 3644 3044 3699
rect 3096 3644 3104 3699
rect 3179 3685 3187 3707
rect 3180 3678 3205 3685
rect 3137 3664 3189 3667
rect 1997 3618 2005 3624
rect 2037 3618 2049 3624
rect 2119 3618 2131 3624
rect 2191 3618 2203 3624
rect 2231 3618 2243 3624
rect 2271 3618 2283 3624
rect 2311 3618 2323 3624
rect 2351 3618 2363 3624
rect 2401 3618 2413 3624
rect 2463 3618 2475 3624
rect 2511 3618 2523 3624
rect 2569 3618 2581 3624
rect 2671 3618 2683 3624
rect 2751 3618 2763 3624
rect 2791 3618 2803 3624
rect 2831 3618 2843 3624
rect 2871 3618 2883 3624
rect 2911 3618 2923 3624
rect 2951 3618 2963 3624
rect 2991 3618 3003 3624
rect 3149 3658 3177 3664
rect 3197 3664 3205 3678
rect 3254 3664 3262 3707
rect 3456 3713 3464 3796
rect 3398 3664 3406 3707
rect 3254 3653 3280 3664
rect 3017 3618 3029 3624
rect 3111 3618 3123 3624
rect 3157 3618 3169 3624
rect 3258 3618 3270 3624
rect 3308 3618 3320 3624
rect 3380 3653 3406 3664
rect 3456 3644 3464 3699
rect 3518 3682 3526 3796
rect 3702 3836 3714 3842
rect 3752 3836 3764 3842
rect 3821 3836 3833 3842
rect 3887 3836 3899 3842
rect 3933 3836 3945 3842
rect 3991 3836 4003 3842
rect 4059 3836 4071 3842
rect 4171 3836 4183 3842
rect 4217 3836 4229 3842
rect 4317 3836 4329 3842
rect 4375 3836 4387 3842
rect 4421 3836 4433 3842
rect 4487 3836 4499 3842
rect 4559 3836 4571 3842
rect 4651 3836 4663 3842
rect 3857 3790 3865 3796
rect 3907 3790 3919 3796
rect 3847 3776 3865 3790
rect 3893 3778 3915 3790
rect 3961 3782 3973 3816
rect 3857 3770 3865 3776
rect 3857 3762 3895 3770
rect 3913 3766 3943 3772
rect 3561 3721 3569 3756
rect 3633 3721 3641 3756
rect 3733 3721 3741 3756
rect 3801 3748 3863 3756
rect 3567 3707 3569 3721
rect 3497 3674 3535 3682
rect 3497 3664 3509 3674
rect 3561 3664 3569 3707
rect 3639 3685 3647 3707
rect 3739 3685 3747 3707
rect 3640 3678 3665 3685
rect 3740 3678 3765 3685
rect 3340 3618 3352 3624
rect 3390 3618 3402 3624
rect 3559 3654 3569 3664
rect 3597 3664 3649 3667
rect 3609 3658 3637 3664
rect 3657 3664 3665 3678
rect 3697 3664 3749 3667
rect 3709 3658 3737 3664
rect 3757 3664 3765 3678
rect 3801 3664 3807 3748
rect 3913 3752 3919 3766
rect 3961 3758 3967 3776
rect 3875 3746 3919 3752
rect 3927 3752 3967 3758
rect 3846 3707 3873 3714
rect 3820 3696 3826 3701
rect 3820 3688 3854 3696
rect 3859 3680 3866 3688
rect 3927 3680 3933 3752
rect 3987 3744 4001 3752
rect 3993 3693 4007 3707
rect 4015 3693 4023 3756
rect 4037 3750 4045 3796
rect 4197 3762 4209 3764
rect 4197 3756 4237 3762
rect 4347 3782 4359 3816
rect 4401 3790 4413 3796
rect 4455 3790 4463 3796
rect 4405 3778 4427 3790
rect 4455 3776 4473 3790
rect 4353 3758 4359 3776
rect 4377 3766 4407 3772
rect 4455 3770 4463 3776
rect 4037 3744 4063 3750
rect 4060 3738 4063 3744
rect 3859 3674 3933 3680
rect 4007 3679 4023 3693
rect 3859 3668 3866 3674
rect 3927 3672 3933 3674
rect 3891 3656 3912 3663
rect 4015 3664 4023 3679
rect 4060 3682 4067 3738
rect 4081 3721 4089 3756
rect 4143 3749 4160 3756
rect 4087 3707 4089 3721
rect 4060 3676 4063 3682
rect 3840 3644 3847 3650
rect 3905 3644 3912 3656
rect 3962 3650 3973 3658
rect 3962 3644 3969 3650
rect 3840 3638 3853 3644
rect 4041 3670 4063 3676
rect 4041 3644 4049 3670
rect 4081 3664 4089 3707
rect 4153 3701 4160 3749
rect 4258 3721 4266 3756
rect 4153 3644 4160 3687
rect 4258 3664 4266 3707
rect 3437 3618 3449 3624
rect 3527 3618 3539 3624
rect 3617 3618 3629 3624
rect 3717 3618 3729 3624
rect 3821 3618 3833 3624
rect 3883 3618 3895 3624
rect 3931 3618 3943 3624
rect 3989 3618 4001 3624
rect 4059 3618 4071 3624
rect 4131 3618 4143 3624
rect 4171 3618 4183 3624
rect 4240 3653 4266 3664
rect 4297 3693 4305 3756
rect 4319 3744 4333 3752
rect 4353 3752 4393 3758
rect 4313 3693 4327 3707
rect 4297 3679 4313 3693
rect 4387 3680 4393 3752
rect 4401 3752 4407 3766
rect 4425 3762 4463 3770
rect 4401 3746 4445 3752
rect 4457 3748 4519 3756
rect 4447 3707 4474 3714
rect 4494 3696 4500 3701
rect 4466 3688 4500 3696
rect 4454 3680 4461 3688
rect 4297 3664 4305 3679
rect 4387 3674 4461 3680
rect 4387 3672 4393 3674
rect 4454 3668 4461 3674
rect 4347 3650 4358 3658
rect 4351 3644 4358 3650
rect 4408 3656 4429 3663
rect 4513 3664 4519 3748
rect 4537 3750 4545 3796
rect 4677 3836 4689 3842
rect 4537 3744 4563 3750
rect 4560 3738 4563 3744
rect 4560 3682 4567 3738
rect 4581 3721 4589 3756
rect 4587 3707 4589 3721
rect 4636 3713 4644 3796
rect 4696 3713 4704 3796
rect 4560 3676 4563 3682
rect 4408 3644 4415 3656
rect 4473 3644 4480 3650
rect 4467 3638 4480 3644
rect 4541 3670 4563 3676
rect 4541 3644 4549 3670
rect 4581 3664 4589 3707
rect 4636 3644 4644 3699
rect 4696 3644 4704 3699
rect 4200 3618 4212 3624
rect 4250 3618 4262 3624
rect 4319 3618 4331 3624
rect 4377 3618 4389 3624
rect 4425 3618 4437 3624
rect 4487 3618 4499 3624
rect 4559 3618 4571 3624
rect 4651 3618 4663 3624
rect 4677 3618 4689 3624
rect 4782 3618 4842 4082
rect 4 3616 4842 3618
rect 4776 3604 4842 3616
rect 4 3602 4842 3604
rect 69 3596 81 3602
rect 121 3596 133 3602
rect 183 3596 195 3602
rect 231 3596 243 3602
rect 289 3596 301 3602
rect 371 3596 383 3602
rect 449 3596 461 3602
rect 531 3596 543 3602
rect 631 3596 643 3602
rect 679 3596 691 3602
rect 777 3596 789 3602
rect 877 3596 889 3602
rect 1010 3596 1022 3602
rect 140 3576 153 3582
rect 140 3570 147 3576
rect 205 3564 212 3576
rect 39 3548 51 3556
rect 39 3542 63 3548
rect 55 3493 63 3542
rect 55 3424 63 3479
rect 101 3472 107 3556
rect 191 3557 212 3564
rect 262 3570 269 3576
rect 262 3562 273 3570
rect 159 3546 166 3552
rect 227 3546 233 3548
rect 159 3540 233 3546
rect 315 3541 323 3556
rect 159 3532 166 3540
rect 120 3524 154 3532
rect 120 3519 126 3524
rect 146 3506 173 3513
rect 101 3464 163 3472
rect 175 3468 219 3474
rect 157 3450 195 3458
rect 213 3454 219 3468
rect 227 3468 233 3540
rect 307 3527 323 3541
rect 293 3513 307 3527
rect 227 3462 267 3468
rect 287 3468 301 3476
rect 315 3464 323 3527
rect 356 3521 364 3576
rect 419 3548 431 3556
rect 419 3542 443 3548
rect 157 3444 165 3450
rect 213 3448 243 3454
rect 261 3444 267 3462
rect 147 3430 165 3444
rect 193 3430 215 3442
rect 157 3424 165 3430
rect 207 3424 219 3430
rect 261 3404 273 3438
rect 356 3424 364 3507
rect 435 3493 443 3542
rect 495 3542 503 3556
rect 523 3556 551 3562
rect 511 3553 563 3556
rect 595 3542 603 3556
rect 623 3556 651 3562
rect 611 3553 663 3556
rect 709 3548 721 3556
rect 769 3556 797 3560
rect 809 3590 837 3596
rect 757 3554 809 3556
rect 697 3542 721 3548
rect 819 3546 825 3556
rect 495 3535 520 3542
rect 595 3535 620 3542
rect 513 3513 521 3535
rect 613 3513 621 3535
rect 435 3424 443 3479
rect 519 3464 527 3499
rect 619 3464 627 3499
rect 697 3493 705 3542
rect 796 3539 825 3546
rect 796 3513 804 3539
rect 896 3521 904 3576
rect 937 3557 953 3563
rect 31 3378 43 3384
rect 71 3378 83 3384
rect 121 3378 133 3384
rect 187 3378 199 3384
rect 233 3378 245 3384
rect 291 3378 303 3384
rect 371 3378 383 3384
rect 411 3378 423 3384
rect 451 3378 463 3384
rect 496 3378 508 3384
rect 546 3378 558 3384
rect 697 3424 705 3479
rect 797 3464 805 3499
rect 596 3378 608 3384
rect 646 3378 658 3384
rect 677 3378 689 3384
rect 717 3378 729 3384
rect 896 3424 904 3507
rect 937 3467 943 3557
rect 956 3538 974 3540
rect 956 3529 986 3538
rect 1040 3596 1052 3602
rect 1090 3596 1102 3602
rect 1137 3596 1149 3602
rect 1177 3596 1189 3602
rect 1219 3596 1231 3602
rect 1299 3596 1311 3602
rect 1397 3596 1409 3602
rect 1501 3596 1513 3602
rect 1563 3596 1575 3602
rect 1611 3596 1623 3602
rect 1669 3596 1681 3602
rect 1769 3596 1781 3602
rect 1817 3596 1829 3602
rect 1897 3596 1909 3602
rect 2009 3596 2021 3602
rect 2081 3596 2093 3602
rect 2139 3596 2151 3602
rect 2218 3596 2230 3602
rect 2317 3596 2329 3602
rect 2377 3596 2389 3602
rect 2459 3596 2471 3602
rect 2517 3596 2529 3602
rect 2565 3596 2577 3602
rect 2627 3596 2639 3602
rect 2697 3596 2709 3602
rect 2799 3596 2811 3602
rect 2859 3596 2871 3602
rect 2959 3596 2971 3602
rect 3017 3596 3029 3602
rect 3065 3596 3077 3602
rect 3127 3596 3139 3602
rect 3231 3596 3243 3602
rect 3311 3596 3323 3602
rect 1080 3556 1106 3567
rect 956 3501 964 3529
rect 1098 3513 1106 3556
rect 1160 3533 1167 3576
rect 1249 3548 1261 3556
rect 1329 3548 1341 3556
rect 1389 3556 1417 3562
rect 1377 3553 1429 3556
rect 1520 3576 1533 3582
rect 1520 3570 1527 3576
rect 1585 3564 1592 3576
rect 955 3432 962 3487
rect 1098 3464 1106 3499
rect 1160 3471 1167 3519
rect 1237 3542 1261 3548
rect 1317 3542 1341 3548
rect 1437 3542 1445 3556
rect 1237 3493 1245 3542
rect 1317 3493 1325 3542
rect 1420 3535 1445 3542
rect 1419 3513 1427 3535
rect 1160 3464 1177 3471
rect 1037 3458 1077 3464
rect 1037 3456 1049 3458
rect 955 3426 1002 3432
rect 955 3424 963 3426
rect 757 3378 769 3384
rect 827 3378 839 3384
rect 991 3424 1002 3426
rect 1237 3424 1245 3479
rect 1317 3424 1325 3479
rect 1413 3464 1421 3499
rect 1481 3472 1487 3556
rect 1571 3557 1592 3564
rect 1642 3570 1649 3576
rect 1642 3562 1653 3570
rect 1539 3546 1546 3552
rect 1607 3546 1613 3548
rect 1539 3540 1613 3546
rect 1695 3541 1703 3556
rect 1809 3556 1837 3562
rect 1739 3548 1751 3556
rect 1797 3553 1849 3556
rect 2051 3556 2061 3566
rect 1739 3542 1763 3548
rect 1857 3542 1865 3556
rect 1539 3532 1546 3540
rect 1500 3524 1534 3532
rect 1500 3519 1506 3524
rect 1526 3506 1553 3513
rect 1481 3464 1543 3472
rect 1555 3468 1599 3474
rect 877 3378 889 3384
rect 971 3378 983 3384
rect 1011 3378 1023 3384
rect 1057 3378 1069 3384
rect 1137 3378 1149 3384
rect 1217 3378 1229 3384
rect 1257 3378 1269 3384
rect 1297 3378 1309 3384
rect 1337 3378 1349 3384
rect 1537 3450 1575 3458
rect 1593 3454 1599 3468
rect 1607 3468 1613 3540
rect 1687 3527 1703 3541
rect 1673 3513 1687 3527
rect 1607 3462 1647 3468
rect 1667 3468 1681 3476
rect 1695 3464 1703 3527
rect 1755 3493 1763 3542
rect 1840 3535 1865 3542
rect 1839 3513 1847 3535
rect 1916 3513 1924 3556
rect 1979 3548 1991 3556
rect 1979 3542 2003 3548
rect 1537 3444 1545 3450
rect 1593 3448 1623 3454
rect 1641 3444 1647 3462
rect 1527 3430 1545 3444
rect 1573 3430 1595 3442
rect 1537 3424 1545 3430
rect 1587 3424 1599 3430
rect 1641 3404 1653 3438
rect 1755 3424 1763 3479
rect 1833 3464 1841 3499
rect 1916 3464 1924 3499
rect 1995 3493 2003 3542
rect 2051 3513 2059 3556
rect 2111 3546 2123 3556
rect 2169 3548 2181 3556
rect 2085 3538 2123 3546
rect 2157 3542 2181 3548
rect 2051 3499 2053 3513
rect 1382 3378 1394 3384
rect 1432 3378 1444 3384
rect 1501 3378 1513 3384
rect 1567 3378 1579 3384
rect 1613 3378 1625 3384
rect 1671 3378 1683 3384
rect 1731 3378 1743 3384
rect 1771 3378 1783 3384
rect 1802 3378 1814 3384
rect 1852 3378 1864 3384
rect 1995 3424 2003 3479
rect 2051 3464 2059 3499
rect 2094 3424 2102 3538
rect 2157 3493 2165 3542
rect 2266 3538 2284 3540
rect 2254 3529 2284 3538
rect 2276 3501 2284 3529
rect 2336 3521 2344 3576
rect 2396 3521 2404 3576
rect 2607 3576 2620 3582
rect 2491 3570 2498 3576
rect 2487 3562 2498 3570
rect 2548 3564 2555 3576
rect 2613 3570 2620 3576
rect 2437 3541 2445 3556
rect 2548 3557 2569 3564
rect 2527 3546 2533 3548
rect 2594 3546 2601 3552
rect 2437 3527 2453 3541
rect 2527 3540 2601 3546
rect 2157 3424 2165 3479
rect 2278 3432 2285 3487
rect 2238 3426 2285 3432
rect 2238 3424 2249 3426
rect 1897 3378 1909 3384
rect 1971 3378 1983 3384
rect 2011 3378 2023 3384
rect 2067 3378 2079 3384
rect 2111 3378 2123 3384
rect 2137 3378 2149 3384
rect 2177 3378 2189 3384
rect 2277 3424 2285 3426
rect 2336 3424 2344 3507
rect 2396 3424 2404 3507
rect 2437 3464 2445 3527
rect 2453 3513 2467 3527
rect 2459 3468 2473 3476
rect 2527 3468 2533 3540
rect 2594 3532 2601 3540
rect 2606 3524 2640 3532
rect 2634 3519 2640 3524
rect 2587 3506 2614 3513
rect 2493 3462 2533 3468
rect 2541 3468 2585 3474
rect 2493 3444 2499 3462
rect 2541 3454 2547 3468
rect 2653 3472 2659 3556
rect 2689 3556 2717 3562
rect 2677 3553 2729 3556
rect 2737 3542 2745 3556
rect 2781 3550 2789 3576
rect 2781 3544 2803 3550
rect 2720 3535 2745 3542
rect 2800 3538 2803 3544
rect 2719 3513 2727 3535
rect 2597 3464 2659 3472
rect 2713 3464 2721 3499
rect 2800 3482 2807 3538
rect 2821 3513 2829 3556
rect 2889 3548 2901 3556
rect 2877 3542 2901 3548
rect 3107 3576 3120 3582
rect 2991 3570 2998 3576
rect 2987 3562 2998 3570
rect 3048 3564 3055 3576
rect 3113 3570 3120 3576
rect 2827 3499 2829 3513
rect 2800 3476 2803 3482
rect 2777 3470 2803 3476
rect 2517 3448 2547 3454
rect 2565 3450 2603 3458
rect 2595 3444 2603 3450
rect 2487 3404 2499 3438
rect 2545 3430 2567 3442
rect 2595 3430 2613 3444
rect 2541 3424 2553 3430
rect 2595 3424 2603 3430
rect 2777 3424 2785 3470
rect 2821 3464 2829 3499
rect 2877 3493 2885 3542
rect 2937 3541 2945 3556
rect 3048 3557 3069 3564
rect 3027 3546 3033 3548
rect 3094 3546 3101 3552
rect 2937 3527 2953 3541
rect 3027 3540 3101 3546
rect 2877 3424 2885 3479
rect 2937 3464 2945 3527
rect 2953 3513 2967 3527
rect 2959 3468 2973 3476
rect 3027 3468 3033 3540
rect 3094 3532 3101 3540
rect 3106 3524 3140 3532
rect 3134 3519 3140 3524
rect 3087 3506 3114 3513
rect 2993 3462 3033 3468
rect 3041 3468 3085 3474
rect 2993 3444 2999 3462
rect 3041 3454 3047 3468
rect 3153 3472 3159 3556
rect 3195 3542 3203 3556
rect 3223 3556 3251 3562
rect 3337 3596 3349 3602
rect 3377 3596 3389 3602
rect 3417 3596 3429 3602
rect 3491 3596 3503 3602
rect 3531 3596 3543 3602
rect 3560 3596 3572 3602
rect 3610 3596 3622 3602
rect 3211 3553 3263 3556
rect 3195 3535 3220 3542
rect 3213 3513 3221 3535
rect 3296 3521 3304 3576
rect 3360 3533 3367 3576
rect 3097 3464 3159 3472
rect 3219 3464 3227 3499
rect 3017 3448 3047 3454
rect 3065 3450 3103 3458
rect 3095 3444 3103 3450
rect 2987 3404 2999 3438
rect 3045 3430 3067 3442
rect 3095 3430 3113 3444
rect 3041 3424 3053 3430
rect 3095 3424 3103 3430
rect 3296 3424 3304 3507
rect 3360 3471 3367 3519
rect 3397 3483 3403 3533
rect 3436 3521 3444 3576
rect 3513 3533 3520 3576
rect 3657 3596 3665 3602
rect 3697 3596 3709 3602
rect 3792 3596 3804 3602
rect 3848 3596 3860 3602
rect 3929 3596 3941 3602
rect 3979 3596 3991 3602
rect 4037 3596 4049 3602
rect 4085 3596 4097 3602
rect 4147 3596 4159 3602
rect 4219 3596 4231 3602
rect 4277 3596 4289 3602
rect 4325 3596 4337 3602
rect 4387 3596 4399 3602
rect 4451 3596 4463 3602
rect 4491 3596 4503 3602
rect 4531 3596 4543 3602
rect 4571 3596 4583 3602
rect 4611 3596 4623 3602
rect 4657 3596 4669 3602
rect 3600 3556 3626 3567
rect 3397 3477 3413 3483
rect 3360 3464 3377 3471
rect 2217 3378 2229 3384
rect 2257 3378 2269 3384
rect 2317 3378 2329 3384
rect 2377 3378 2389 3384
rect 2457 3378 2469 3384
rect 2515 3378 2527 3384
rect 2561 3378 2573 3384
rect 2627 3378 2639 3384
rect 2682 3378 2694 3384
rect 2732 3378 2744 3384
rect 2799 3378 2811 3384
rect 2857 3378 2869 3384
rect 2897 3378 2909 3384
rect 2957 3378 2969 3384
rect 3015 3378 3027 3384
rect 3061 3378 3073 3384
rect 3127 3378 3139 3384
rect 3196 3378 3208 3384
rect 3246 3378 3258 3384
rect 3311 3378 3323 3384
rect 3436 3424 3444 3507
rect 3513 3471 3520 3519
rect 3618 3513 3626 3556
rect 3683 3548 3689 3576
rect 4127 3576 4140 3582
rect 4011 3570 4018 3576
rect 4007 3562 4018 3570
rect 4068 3564 4075 3576
rect 4133 3570 4140 3576
rect 3683 3542 3693 3548
rect 3503 3464 3520 3471
rect 3618 3464 3626 3499
rect 3698 3481 3704 3536
rect 3720 3521 3727 3556
rect 3657 3472 3693 3480
rect 3657 3464 3665 3472
rect 3557 3458 3597 3464
rect 3557 3456 3569 3458
rect 3714 3463 3723 3507
rect 3820 3513 3827 3556
rect 3899 3548 3911 3556
rect 3899 3542 3923 3548
rect 3813 3476 3819 3499
rect 3915 3493 3923 3542
rect 3957 3541 3965 3556
rect 4068 3557 4089 3564
rect 4047 3546 4053 3548
rect 4114 3546 4121 3552
rect 3957 3527 3973 3541
rect 4047 3540 4121 3546
rect 3792 3470 3819 3476
rect 3792 3464 3804 3470
rect 3719 3454 3723 3463
rect 3783 3384 3811 3390
rect 3823 3456 3851 3462
rect 3915 3424 3923 3479
rect 3957 3464 3965 3527
rect 3973 3513 3987 3527
rect 3979 3468 3993 3476
rect 4047 3468 4053 3540
rect 4114 3532 4121 3540
rect 4126 3524 4160 3532
rect 4154 3519 4160 3524
rect 4107 3506 4134 3513
rect 4013 3462 4053 3468
rect 4061 3468 4105 3474
rect 4013 3444 4019 3462
rect 4061 3454 4067 3468
rect 4173 3472 4179 3556
rect 4117 3464 4179 3472
rect 4037 3448 4067 3454
rect 4085 3450 4123 3458
rect 4115 3444 4123 3450
rect 4007 3404 4019 3438
rect 4065 3430 4087 3442
rect 4115 3430 4133 3444
rect 4061 3424 4073 3430
rect 4115 3424 4123 3430
rect 4367 3576 4380 3582
rect 4251 3570 4258 3576
rect 4247 3562 4258 3570
rect 4308 3564 4315 3576
rect 4373 3570 4380 3576
rect 4197 3541 4205 3556
rect 4308 3557 4329 3564
rect 4649 3556 4677 3562
rect 4287 3546 4293 3548
rect 4354 3546 4361 3552
rect 4197 3527 4213 3541
rect 4287 3540 4361 3546
rect 4197 3464 4205 3527
rect 4213 3513 4227 3527
rect 4219 3468 4233 3476
rect 4287 3468 4293 3540
rect 4354 3532 4361 3540
rect 4366 3524 4400 3532
rect 4394 3519 4400 3524
rect 4347 3506 4374 3513
rect 4253 3462 4293 3468
rect 4301 3468 4345 3474
rect 4253 3444 4259 3462
rect 4301 3454 4307 3468
rect 4413 3472 4419 3556
rect 4472 3550 4484 3556
rect 4512 3550 4524 3556
rect 4551 3550 4563 3556
rect 4592 3550 4604 3556
rect 4637 3553 4689 3556
rect 4466 3549 4484 3550
rect 4465 3542 4484 3549
rect 4498 3542 4524 3550
rect 4538 3542 4563 3550
rect 4577 3542 4604 3550
rect 4697 3542 4705 3556
rect 4465 3521 4472 3542
rect 4498 3536 4506 3542
rect 4538 3536 4546 3542
rect 4577 3536 4585 3542
rect 4490 3524 4506 3536
rect 4530 3524 4546 3536
rect 4570 3524 4585 3536
rect 4680 3535 4705 3542
rect 4467 3507 4472 3521
rect 4357 3464 4419 3472
rect 4465 3478 4472 3507
rect 4498 3478 4506 3524
rect 4538 3478 4546 3524
rect 4577 3478 4585 3524
rect 4679 3513 4687 3535
rect 4465 3470 4483 3478
rect 4498 3470 4523 3478
rect 4538 3470 4563 3478
rect 4577 3470 4603 3478
rect 4471 3464 4483 3470
rect 4511 3464 4523 3470
rect 4551 3464 4563 3470
rect 4591 3464 4603 3470
rect 4673 3464 4681 3499
rect 4277 3448 4307 3454
rect 4325 3450 4363 3458
rect 4355 3444 4363 3450
rect 4247 3404 4259 3438
rect 4305 3430 4327 3442
rect 4355 3430 4373 3444
rect 4301 3424 4313 3430
rect 4355 3424 4363 3430
rect 3337 3378 3349 3384
rect 3417 3378 3429 3384
rect 3531 3378 3543 3384
rect 3577 3378 3589 3384
rect 3687 3378 3699 3384
rect 3831 3378 3843 3384
rect 3891 3378 3903 3384
rect 3931 3378 3943 3384
rect 3977 3378 3989 3384
rect 4035 3378 4047 3384
rect 4081 3378 4093 3384
rect 4147 3378 4159 3384
rect 4217 3378 4229 3384
rect 4275 3378 4287 3384
rect 4321 3378 4333 3384
rect 4387 3378 4399 3384
rect 4451 3378 4463 3384
rect 4491 3378 4503 3384
rect 4531 3378 4543 3384
rect 4571 3378 4583 3384
rect 4611 3378 4623 3384
rect 4642 3378 4654 3384
rect 4692 3378 4704 3384
rect -62 3376 4776 3378
rect -62 3364 4 3376
rect -62 3362 4776 3364
rect -62 2898 -2 3362
rect 41 3356 53 3362
rect 107 3356 119 3362
rect 153 3356 165 3362
rect 211 3356 223 3362
rect 331 3356 343 3362
rect 391 3356 403 3362
rect 431 3356 443 3362
rect 477 3356 489 3362
rect 535 3356 547 3362
rect 581 3356 593 3362
rect 647 3356 659 3362
rect 716 3356 728 3362
rect 766 3356 778 3362
rect 871 3356 883 3362
rect 917 3356 929 3362
rect 957 3356 969 3362
rect 1031 3356 1043 3362
rect 1071 3356 1083 3362
rect 1127 3356 1139 3362
rect 1171 3356 1183 3362
rect 77 3310 85 3316
rect 127 3310 139 3316
rect 67 3296 85 3310
rect 113 3298 135 3310
rect 181 3302 193 3336
rect 77 3290 85 3296
rect 77 3282 115 3290
rect 133 3286 163 3292
rect 21 3268 83 3276
rect 21 3184 27 3268
rect 133 3272 139 3286
rect 181 3278 187 3296
rect 95 3266 139 3272
rect 147 3272 187 3278
rect 66 3227 93 3234
rect 40 3216 46 3221
rect 40 3208 74 3216
rect 79 3200 86 3208
rect 147 3200 153 3272
rect 283 3350 311 3356
rect 323 3278 351 3284
rect 397 3283 403 3293
rect 377 3277 403 3283
rect 207 3264 221 3272
rect 213 3213 227 3227
rect 235 3213 243 3276
rect 292 3270 304 3276
rect 292 3264 319 3270
rect 313 3241 319 3264
rect 79 3194 153 3200
rect 227 3199 243 3213
rect 79 3188 86 3194
rect 147 3192 153 3194
rect 111 3176 132 3183
rect 235 3184 243 3199
rect 320 3184 327 3227
rect 377 3227 383 3277
rect 415 3261 423 3316
rect 507 3302 519 3336
rect 561 3310 573 3316
rect 615 3310 623 3316
rect 565 3298 587 3310
rect 615 3296 633 3310
rect 513 3278 519 3296
rect 537 3286 567 3292
rect 615 3290 623 3296
rect 415 3198 423 3247
rect 399 3192 423 3198
rect 457 3213 465 3276
rect 479 3264 493 3272
rect 513 3272 553 3278
rect 473 3213 487 3227
rect 457 3199 473 3213
rect 547 3200 553 3272
rect 561 3272 567 3286
rect 585 3282 623 3290
rect 823 3350 851 3356
rect 863 3278 891 3284
rect 561 3266 605 3272
rect 617 3268 679 3276
rect 607 3227 634 3234
rect 654 3216 660 3221
rect 626 3208 660 3216
rect 614 3200 621 3208
rect 399 3184 411 3192
rect 457 3184 465 3199
rect 547 3194 621 3200
rect 547 3192 553 3194
rect 60 3164 67 3170
rect 125 3164 132 3176
rect 182 3170 193 3178
rect 182 3164 189 3170
rect 60 3158 73 3164
rect 614 3188 621 3194
rect 507 3170 518 3178
rect 511 3164 518 3170
rect 568 3176 589 3183
rect 673 3184 679 3268
rect 739 3241 747 3276
rect 832 3270 844 3276
rect 832 3264 859 3270
rect 853 3241 859 3264
rect 937 3261 945 3316
rect 1015 3314 1023 3316
rect 1051 3314 1062 3316
rect 1015 3308 1062 3314
rect 733 3205 741 3227
rect 715 3198 740 3205
rect 715 3184 723 3198
rect 568 3164 575 3176
rect 633 3164 640 3170
rect 627 3158 640 3164
rect 731 3184 783 3187
rect 860 3184 867 3227
rect 1015 3253 1022 3308
rect 1197 3356 1209 3362
rect 1237 3356 1249 3362
rect 1302 3356 1314 3362
rect 1352 3356 1364 3362
rect 937 3198 945 3247
rect 1111 3241 1119 3276
rect 1016 3211 1024 3239
rect 1111 3227 1113 3241
rect 1016 3202 1046 3211
rect 1016 3200 1034 3202
rect 937 3192 961 3198
rect 949 3184 961 3192
rect 743 3178 771 3184
rect 41 3138 53 3144
rect 103 3138 115 3144
rect 151 3138 163 3144
rect 209 3138 221 3144
rect 292 3138 304 3144
rect 348 3138 360 3144
rect 429 3138 441 3144
rect 479 3138 491 3144
rect 537 3138 549 3144
rect 585 3138 597 3144
rect 647 3138 659 3144
rect 751 3138 763 3144
rect 832 3138 844 3144
rect 888 3138 900 3144
rect 1111 3184 1119 3227
rect 1154 3202 1162 3316
rect 1218 3314 1229 3316
rect 1257 3314 1265 3316
rect 1218 3308 1265 3314
rect 1258 3253 1265 3308
rect 1397 3356 1409 3362
rect 1437 3356 1449 3362
rect 1521 3356 1533 3362
rect 1591 3356 1603 3362
rect 1631 3356 1643 3362
rect 1333 3241 1341 3276
rect 1417 3261 1425 3316
rect 1497 3277 1501 3286
rect 1256 3211 1264 3239
rect 1145 3194 1183 3202
rect 1171 3184 1183 3194
rect 1111 3174 1121 3184
rect 1234 3202 1264 3211
rect 1339 3205 1347 3227
rect 1246 3200 1264 3202
rect 1340 3198 1365 3205
rect 1297 3184 1349 3187
rect 1309 3178 1337 3184
rect 1357 3184 1365 3198
rect 1417 3198 1425 3247
rect 1497 3233 1506 3277
rect 1662 3356 1674 3362
rect 1712 3356 1724 3362
rect 1555 3268 1563 3276
rect 1527 3260 1563 3268
rect 1577 3277 1593 3283
rect 1417 3192 1441 3198
rect 1429 3184 1441 3192
rect 1493 3184 1500 3219
rect 1516 3204 1522 3259
rect 1527 3192 1537 3198
rect 1531 3164 1537 3192
rect 1577 3183 1583 3277
rect 1615 3261 1623 3316
rect 1776 3356 1788 3362
rect 1826 3356 1838 3362
rect 1727 3297 1773 3303
rect 1857 3356 1869 3362
rect 1897 3356 1909 3362
rect 1942 3356 1954 3362
rect 1992 3356 2004 3362
rect 1615 3198 1623 3247
rect 1693 3241 1701 3276
rect 1799 3241 1807 3276
rect 1877 3261 1885 3316
rect 1907 3277 1923 3283
rect 1699 3205 1707 3227
rect 1793 3205 1801 3227
rect 1700 3198 1725 3205
rect 1567 3177 1583 3183
rect 1599 3192 1623 3198
rect 1599 3184 1611 3192
rect 1657 3184 1709 3187
rect 1669 3178 1697 3184
rect 1717 3184 1725 3198
rect 1775 3198 1800 3205
rect 1877 3198 1885 3247
rect 1917 3203 1923 3277
rect 2056 3356 2068 3362
rect 2106 3356 2118 3362
rect 2137 3356 2149 3362
rect 2202 3356 2214 3362
rect 2252 3356 2264 3362
rect 2331 3356 2343 3362
rect 1973 3241 1981 3276
rect 2079 3241 2087 3276
rect 1775 3184 1783 3198
rect 1877 3192 1901 3198
rect 1917 3197 1933 3203
rect 1979 3205 1987 3227
rect 2073 3205 2081 3227
rect 2156 3233 2164 3316
rect 2357 3356 2369 3362
rect 2397 3356 2409 3362
rect 2457 3356 2469 3362
rect 2515 3356 2527 3362
rect 2561 3356 2573 3362
rect 2627 3356 2639 3362
rect 2699 3356 2711 3362
rect 2777 3356 2789 3362
rect 2835 3356 2847 3362
rect 2881 3356 2893 3362
rect 2947 3356 2959 3362
rect 3016 3356 3028 3362
rect 3066 3356 3078 3362
rect 2233 3241 2241 3276
rect 2316 3233 2324 3316
rect 2377 3261 2385 3316
rect 2487 3302 2499 3336
rect 2541 3310 2553 3316
rect 2595 3310 2603 3316
rect 2545 3298 2567 3310
rect 2595 3296 2613 3310
rect 2493 3278 2499 3296
rect 2517 3286 2547 3292
rect 2595 3290 2603 3296
rect 1980 3198 2005 3205
rect 1791 3184 1843 3187
rect 1889 3184 1901 3192
rect 1803 3178 1831 3184
rect 1937 3184 1989 3187
rect 1949 3178 1977 3184
rect 1997 3184 2005 3198
rect 2055 3198 2080 3205
rect 2055 3184 2063 3198
rect 2071 3184 2123 3187
rect 2083 3178 2111 3184
rect 2156 3164 2164 3219
rect 2239 3205 2247 3227
rect 2240 3198 2265 3205
rect 2197 3184 2249 3187
rect 2209 3178 2237 3184
rect 2257 3184 2265 3198
rect 2316 3164 2324 3219
rect 2377 3198 2385 3247
rect 2437 3213 2445 3276
rect 2459 3264 2473 3272
rect 2493 3272 2533 3278
rect 2453 3213 2467 3227
rect 2437 3199 2453 3213
rect 2527 3200 2533 3272
rect 2541 3272 2547 3286
rect 2565 3282 2603 3290
rect 2541 3266 2585 3272
rect 2597 3268 2659 3276
rect 2587 3227 2614 3234
rect 2634 3216 2640 3221
rect 2606 3208 2640 3216
rect 2594 3200 2601 3208
rect 2377 3192 2401 3198
rect 2389 3184 2401 3192
rect 919 3138 931 3144
rect 1070 3138 1082 3144
rect 1141 3138 1153 3144
rect 1198 3138 1210 3144
rect 1317 3138 1329 3144
rect 1399 3138 1411 3144
rect 1511 3138 1523 3144
rect 1555 3138 1563 3144
rect 1629 3138 1641 3144
rect 1677 3138 1689 3144
rect 1811 3138 1823 3144
rect 1859 3138 1871 3144
rect 1957 3138 1969 3144
rect 2091 3138 2103 3144
rect 2137 3138 2149 3144
rect 2217 3138 2229 3144
rect 2331 3138 2343 3144
rect 2437 3184 2445 3199
rect 2527 3194 2601 3200
rect 2527 3192 2533 3194
rect 2594 3188 2601 3194
rect 2487 3170 2498 3178
rect 2491 3164 2498 3170
rect 2548 3176 2569 3183
rect 2653 3184 2659 3268
rect 2677 3270 2685 3316
rect 2807 3302 2819 3336
rect 2861 3310 2873 3316
rect 2915 3310 2923 3316
rect 2865 3298 2887 3310
rect 2915 3296 2933 3310
rect 2813 3278 2819 3296
rect 2837 3286 2867 3292
rect 2915 3290 2923 3296
rect 2677 3264 2703 3270
rect 2700 3258 2703 3264
rect 2700 3202 2707 3258
rect 2721 3241 2729 3276
rect 2727 3227 2729 3241
rect 2700 3196 2703 3202
rect 2548 3164 2555 3176
rect 2613 3164 2620 3170
rect 2607 3158 2620 3164
rect 2681 3190 2703 3196
rect 2681 3164 2689 3190
rect 2721 3184 2729 3227
rect 2757 3213 2765 3276
rect 2779 3264 2793 3272
rect 2813 3272 2853 3278
rect 2773 3213 2787 3227
rect 2757 3199 2773 3213
rect 2847 3200 2853 3272
rect 2861 3272 2867 3286
rect 2885 3282 2923 3290
rect 3116 3356 3128 3362
rect 3166 3356 3178 3362
rect 3202 3356 3214 3362
rect 3252 3356 3264 3362
rect 3316 3356 3328 3362
rect 3366 3356 3378 3362
rect 3402 3356 3414 3362
rect 3452 3356 3464 3362
rect 3497 3356 3509 3362
rect 3537 3356 3549 3362
rect 3577 3356 3589 3362
rect 3617 3356 3629 3362
rect 3657 3356 3669 3362
rect 3697 3356 3709 3362
rect 3737 3356 3749 3362
rect 3777 3356 3789 3362
rect 3839 3356 3851 3362
rect 3911 3356 3923 3362
rect 3951 3356 3963 3362
rect 4031 3356 4043 3362
rect 4079 3356 4091 3362
rect 4171 3356 4183 3362
rect 2861 3266 2905 3272
rect 2917 3268 2979 3276
rect 2907 3227 2934 3234
rect 2954 3216 2960 3221
rect 2926 3208 2960 3216
rect 2914 3200 2921 3208
rect 2757 3184 2765 3199
rect 2847 3194 2921 3200
rect 2847 3192 2853 3194
rect 2914 3188 2921 3194
rect 2807 3170 2818 3178
rect 2811 3164 2818 3170
rect 2868 3176 2889 3183
rect 2973 3184 2979 3268
rect 3039 3241 3047 3276
rect 3139 3241 3147 3276
rect 3233 3241 3241 3276
rect 3339 3241 3347 3276
rect 3433 3241 3441 3276
rect 3517 3261 3525 3316
rect 3597 3261 3605 3316
rect 3677 3261 3685 3316
rect 3757 3261 3765 3316
rect 3817 3270 3825 3316
rect 3817 3264 3843 3270
rect 3033 3205 3041 3227
rect 3133 3205 3141 3227
rect 3239 3205 3247 3227
rect 3333 3205 3341 3227
rect 3439 3205 3447 3227
rect 3015 3198 3040 3205
rect 3115 3198 3140 3205
rect 3240 3198 3265 3205
rect 3015 3184 3023 3198
rect 2868 3164 2875 3176
rect 2933 3164 2940 3170
rect 2927 3158 2940 3164
rect 3031 3184 3083 3187
rect 3115 3184 3123 3198
rect 3043 3178 3071 3184
rect 3131 3184 3183 3187
rect 3143 3178 3171 3184
rect 3197 3184 3249 3187
rect 3209 3178 3237 3184
rect 3257 3184 3265 3198
rect 3315 3198 3340 3205
rect 3440 3198 3465 3205
rect 3315 3184 3323 3198
rect 3331 3184 3383 3187
rect 3343 3178 3371 3184
rect 3397 3184 3449 3187
rect 3409 3178 3437 3184
rect 3457 3184 3465 3198
rect 3517 3198 3525 3247
rect 3597 3198 3605 3247
rect 3677 3198 3685 3247
rect 3840 3258 3843 3264
rect 3757 3198 3765 3247
rect 3840 3202 3847 3258
rect 3861 3241 3869 3276
rect 3935 3261 3943 3316
rect 4003 3269 4020 3276
rect 3867 3227 3869 3241
rect 3517 3192 3541 3198
rect 3597 3192 3621 3198
rect 3677 3192 3701 3198
rect 3757 3192 3781 3198
rect 3840 3196 3843 3202
rect 3529 3184 3541 3192
rect 3609 3184 3621 3192
rect 3689 3184 3701 3192
rect 3769 3184 3781 3192
rect 3821 3190 3843 3196
rect 3821 3164 3829 3190
rect 3861 3184 3869 3227
rect 3935 3198 3943 3247
rect 3919 3192 3943 3198
rect 4013 3221 4020 3269
rect 4057 3270 4065 3316
rect 4216 3356 4228 3362
rect 4266 3356 4278 3362
rect 4331 3356 4343 3362
rect 4057 3264 4083 3270
rect 4080 3258 4083 3264
rect 3919 3184 3931 3192
rect 4013 3164 4020 3207
rect 4080 3202 4087 3258
rect 4101 3241 4109 3276
rect 4107 3227 4109 3241
rect 4156 3233 4164 3316
rect 4362 3356 4374 3362
rect 4412 3356 4424 3362
rect 4239 3241 4247 3276
rect 4080 3196 4083 3202
rect 4061 3190 4083 3196
rect 4061 3164 4069 3190
rect 4101 3184 4109 3227
rect 2359 3138 2371 3144
rect 2459 3138 2471 3144
rect 2517 3138 2529 3144
rect 2565 3138 2577 3144
rect 2627 3138 2639 3144
rect 2699 3138 2711 3144
rect 2779 3138 2791 3144
rect 2837 3138 2849 3144
rect 2885 3138 2897 3144
rect 2947 3138 2959 3144
rect 3051 3138 3063 3144
rect 3151 3138 3163 3144
rect 3217 3138 3229 3144
rect 3351 3138 3363 3144
rect 3417 3138 3429 3144
rect 3499 3138 3511 3144
rect 3579 3138 3591 3144
rect 3659 3138 3671 3144
rect 3739 3138 3751 3144
rect 3839 3138 3851 3144
rect 3949 3138 3961 3144
rect 4156 3164 4164 3219
rect 4233 3205 4241 3227
rect 4316 3233 4324 3316
rect 4471 3356 4483 3362
rect 4511 3356 4523 3362
rect 4561 3356 4573 3362
rect 4627 3356 4639 3362
rect 4673 3356 4685 3362
rect 4731 3356 4743 3362
rect 4393 3241 4401 3276
rect 4495 3261 4503 3316
rect 4597 3310 4605 3316
rect 4647 3310 4659 3316
rect 4587 3296 4605 3310
rect 4633 3298 4655 3310
rect 4701 3302 4713 3336
rect 4597 3290 4605 3296
rect 4597 3282 4635 3290
rect 4653 3286 4683 3292
rect 4541 3268 4603 3276
rect 4215 3198 4240 3205
rect 4215 3184 4223 3198
rect 4231 3184 4283 3187
rect 4243 3178 4271 3184
rect 4316 3164 4324 3219
rect 4399 3205 4407 3227
rect 4400 3198 4425 3205
rect 4495 3198 4503 3247
rect 4357 3184 4409 3187
rect 4369 3178 4397 3184
rect 4417 3184 4425 3198
rect 4479 3192 4503 3198
rect 4479 3184 4491 3192
rect 4541 3184 4547 3268
rect 4653 3272 4659 3286
rect 4701 3278 4707 3296
rect 4615 3266 4659 3272
rect 4667 3272 4707 3278
rect 4586 3227 4613 3234
rect 4560 3216 4566 3221
rect 4560 3208 4594 3216
rect 4599 3200 4606 3208
rect 4667 3200 4673 3272
rect 4727 3264 4741 3272
rect 4733 3213 4747 3227
rect 4755 3213 4763 3276
rect 4599 3194 4673 3200
rect 4747 3199 4763 3213
rect 4599 3188 4606 3194
rect 4667 3192 4673 3194
rect 4631 3176 4652 3183
rect 4755 3184 4763 3199
rect 4580 3164 4587 3170
rect 4645 3164 4652 3176
rect 4702 3170 4713 3178
rect 4702 3164 4709 3170
rect 4580 3158 4593 3164
rect 3991 3138 4003 3144
rect 4031 3138 4043 3144
rect 4079 3138 4091 3144
rect 4171 3138 4183 3144
rect 4251 3138 4263 3144
rect 4331 3138 4343 3144
rect 4377 3138 4389 3144
rect 4509 3138 4521 3144
rect 4561 3138 4573 3144
rect 4623 3138 4635 3144
rect 4671 3138 4683 3144
rect 4729 3138 4741 3144
rect 4782 3138 4842 3602
rect 4 3136 4842 3138
rect 4776 3124 4842 3136
rect 4 3122 4842 3124
rect 52 3116 64 3122
rect 108 3116 120 3122
rect 181 3116 193 3122
rect 259 3116 271 3122
rect 317 3116 329 3122
rect 365 3116 377 3122
rect 427 3116 439 3122
rect 497 3116 509 3122
rect 579 3116 591 3122
rect 709 3116 721 3122
rect 151 3076 161 3086
rect 80 3033 87 3076
rect 151 3033 159 3076
rect 211 3066 223 3076
rect 185 3058 223 3066
rect 407 3096 420 3102
rect 291 3090 298 3096
rect 287 3082 298 3090
rect 348 3084 355 3096
rect 413 3090 420 3096
rect 237 3061 245 3076
rect 348 3077 369 3084
rect 327 3066 333 3068
rect 394 3066 401 3072
rect 151 3019 153 3033
rect 73 2996 79 3019
rect 52 2990 79 2996
rect 52 2984 64 2990
rect 151 2984 159 3019
rect 43 2904 71 2910
rect 83 2976 111 2982
rect 194 2944 202 3058
rect 237 3047 253 3061
rect 327 3060 401 3066
rect 237 2984 245 3047
rect 253 3033 267 3047
rect 259 2988 273 2996
rect 327 2988 333 3060
rect 394 3052 401 3060
rect 406 3044 440 3052
rect 434 3039 440 3044
rect 387 3026 414 3033
rect 293 2982 333 2988
rect 341 2988 385 2994
rect 293 2964 299 2982
rect 341 2974 347 2988
rect 453 2992 459 3076
rect 489 3076 517 3082
rect 477 3073 529 3076
rect 537 3062 545 3076
rect 609 3068 621 3076
rect 520 3055 545 3062
rect 557 3057 573 3063
rect 519 3033 527 3055
rect 397 2984 459 2992
rect 513 2984 521 3019
rect 317 2968 347 2974
rect 365 2970 403 2978
rect 395 2964 403 2970
rect 287 2924 299 2958
rect 345 2950 367 2962
rect 395 2950 413 2964
rect 341 2944 353 2950
rect 395 2944 403 2950
rect 557 2963 563 3057
rect 597 3062 621 3068
rect 751 3116 763 3122
rect 791 3116 803 3122
rect 819 3116 831 3122
rect 951 3116 963 3122
rect 1051 3116 1063 3122
rect 1111 3116 1123 3122
rect 1151 3116 1163 3122
rect 1231 3116 1243 3122
rect 1279 3116 1291 3122
rect 1391 3116 1403 3122
rect 679 3068 691 3076
rect 679 3062 703 3068
rect 597 3013 605 3062
rect 695 3013 703 3062
rect 773 3053 780 3096
rect 849 3068 861 3076
rect 837 3062 861 3068
rect 915 3062 923 3076
rect 943 3076 971 3082
rect 931 3073 983 3076
rect 1015 3062 1023 3076
rect 1043 3076 1071 3082
rect 1031 3073 1083 3076
rect 547 2957 563 2963
rect 597 2944 605 2999
rect 695 2944 703 2999
rect 773 2991 780 3039
rect 837 3013 845 3062
rect 915 3055 940 3062
rect 1015 3055 1040 3062
rect 933 3033 941 3055
rect 1033 3033 1041 3055
rect 1133 3053 1140 3096
rect 1195 3062 1203 3076
rect 1223 3076 1251 3082
rect 1419 3116 1431 3122
rect 1499 3116 1511 3122
rect 1599 3116 1611 3122
rect 1677 3116 1689 3122
rect 1777 3116 1789 3122
rect 1857 3116 1869 3122
rect 1897 3116 1909 3122
rect 1211 3073 1263 3076
rect 1309 3068 1321 3076
rect 1297 3062 1321 3068
rect 1195 3055 1220 3062
rect 763 2984 780 2991
rect 91 2898 103 2904
rect 167 2898 179 2904
rect 211 2898 223 2904
rect 257 2898 269 2904
rect 315 2898 327 2904
rect 361 2898 373 2904
rect 427 2898 439 2904
rect 482 2898 494 2904
rect 532 2898 544 2904
rect 577 2898 589 2904
rect 617 2898 629 2904
rect 837 2944 845 2999
rect 939 2984 947 3019
rect 1039 2984 1047 3019
rect 1133 2991 1140 3039
rect 1213 3033 1221 3055
rect 1123 2984 1140 2991
rect 1219 2984 1227 3019
rect 1297 3013 1305 3062
rect 1376 3033 1384 3076
rect 1449 3068 1461 3076
rect 1529 3068 1541 3076
rect 1437 3062 1461 3068
rect 1517 3062 1541 3068
rect 1581 3070 1589 3096
rect 1669 3076 1697 3082
rect 1581 3064 1603 3070
rect 671 2898 683 2904
rect 711 2898 723 2904
rect 791 2898 803 2904
rect 817 2898 829 2904
rect 857 2898 869 2904
rect 916 2898 928 2904
rect 966 2898 978 2904
rect 1016 2898 1028 2904
rect 1066 2898 1078 2904
rect 1151 2898 1163 2904
rect 1297 2944 1305 2999
rect 1376 2984 1384 3019
rect 1437 3013 1445 3062
rect 1517 3013 1525 3062
rect 1600 3058 1603 3064
rect 1600 3002 1607 3058
rect 1621 3033 1629 3076
rect 1657 3073 1709 3076
rect 1769 3076 1797 3082
rect 1717 3062 1725 3076
rect 1757 3073 1809 3076
rect 1940 3116 1952 3122
rect 1990 3116 2002 3122
rect 1817 3062 1825 3076
rect 1700 3055 1725 3062
rect 1800 3055 1825 3062
rect 1627 3019 1629 3033
rect 1699 3033 1707 3055
rect 1799 3033 1807 3055
rect 1880 3053 1887 3096
rect 2037 3116 2049 3122
rect 2117 3116 2129 3122
rect 2197 3116 2209 3122
rect 2237 3116 2249 3122
rect 2329 3116 2341 3122
rect 2377 3116 2389 3122
rect 2457 3116 2469 3122
rect 2537 3116 2549 3122
rect 2639 3116 2651 3122
rect 2699 3116 2711 3122
rect 2801 3116 2813 3122
rect 2863 3116 2875 3122
rect 2911 3116 2923 3122
rect 2969 3116 2981 3122
rect 3031 3116 3043 3122
rect 3071 3116 3083 3122
rect 1980 3076 2006 3087
rect 1827 3037 1843 3043
rect 1196 2898 1208 2904
rect 1246 2898 1258 2904
rect 1437 2944 1445 2999
rect 1517 2944 1525 2999
rect 1600 2996 1603 3002
rect 1577 2990 1603 2996
rect 1577 2944 1585 2990
rect 1621 2984 1629 3019
rect 1693 2984 1701 3019
rect 1793 2984 1801 3019
rect 1837 2987 1843 3037
rect 1880 2991 1887 3039
rect 1998 3033 2006 3076
rect 2056 3041 2064 3096
rect 2109 3076 2137 3082
rect 2097 3073 2149 3076
rect 2157 3062 2165 3076
rect 2140 3055 2165 3062
rect 1277 2898 1289 2904
rect 1317 2898 1329 2904
rect 1391 2898 1403 2904
rect 1417 2898 1429 2904
rect 1457 2898 1469 2904
rect 1497 2898 1509 2904
rect 1537 2898 1549 2904
rect 1599 2898 1611 2904
rect 1662 2898 1674 2904
rect 1712 2898 1724 2904
rect 1880 2984 1897 2991
rect 1998 2984 2006 3019
rect 1762 2898 1774 2904
rect 1812 2898 1824 2904
rect 1937 2978 1977 2984
rect 1937 2976 1949 2978
rect 2056 2944 2064 3027
rect 2139 3033 2147 3055
rect 2220 3053 2227 3096
rect 2369 3076 2397 3082
rect 2299 3068 2311 3076
rect 2357 3073 2409 3076
rect 2299 3062 2323 3068
rect 2417 3062 2425 3076
rect 2133 2984 2141 3019
rect 2220 2991 2227 3039
rect 2315 3013 2323 3062
rect 2400 3055 2425 3062
rect 2399 3033 2407 3055
rect 2476 3041 2484 3096
rect 2529 3076 2557 3082
rect 2517 3073 2569 3076
rect 2577 3062 2585 3076
rect 2621 3070 2629 3096
rect 2621 3064 2643 3070
rect 2560 3055 2585 3062
rect 2640 3058 2643 3064
rect 2220 2984 2237 2991
rect 1857 2898 1869 2904
rect 1957 2898 1969 2904
rect 2037 2898 2049 2904
rect 2102 2898 2114 2904
rect 2152 2898 2164 2904
rect 2315 2944 2323 2999
rect 2393 2984 2401 3019
rect 2197 2898 2209 2904
rect 2291 2898 2303 2904
rect 2331 2898 2343 2904
rect 2476 2944 2484 3027
rect 2559 3033 2567 3055
rect 2553 2984 2561 3019
rect 2640 3002 2647 3058
rect 2661 3033 2669 3076
rect 2729 3068 2741 3076
rect 2717 3062 2741 3068
rect 2820 3096 2833 3102
rect 2820 3090 2827 3096
rect 2885 3084 2892 3096
rect 2667 3019 2669 3033
rect 2640 2996 2643 3002
rect 2617 2990 2643 2996
rect 2362 2898 2374 2904
rect 2412 2898 2424 2904
rect 2617 2944 2625 2990
rect 2661 2984 2669 3019
rect 2717 3013 2725 3062
rect 2717 2944 2725 2999
rect 2781 2992 2787 3076
rect 2871 3077 2892 3084
rect 2942 3090 2949 3096
rect 2942 3082 2953 3090
rect 2839 3066 2846 3072
rect 3118 3116 3130 3122
rect 3168 3116 3180 3122
rect 2907 3066 2913 3068
rect 2839 3060 2913 3066
rect 2995 3061 3003 3076
rect 2839 3052 2846 3060
rect 2800 3044 2834 3052
rect 2800 3039 2806 3044
rect 2826 3026 2853 3033
rect 2781 2984 2843 2992
rect 2855 2988 2899 2994
rect 2837 2970 2875 2978
rect 2893 2974 2899 2988
rect 2907 2988 2913 3060
rect 2987 3047 3003 3061
rect 2973 3033 2987 3047
rect 2907 2982 2947 2988
rect 2967 2988 2981 2996
rect 2995 2984 3003 3047
rect 3053 3053 3060 3096
rect 3114 3076 3140 3087
rect 3197 3116 3209 3122
rect 3237 3116 3249 3122
rect 3301 3116 3313 3122
rect 3363 3116 3375 3122
rect 3411 3116 3423 3122
rect 3469 3116 3481 3122
rect 3541 3116 3553 3122
rect 3603 3116 3615 3122
rect 3651 3116 3663 3122
rect 3709 3116 3721 3122
rect 3757 3116 3769 3122
rect 3797 3116 3809 3122
rect 3891 3116 3903 3122
rect 3991 3116 4003 3122
rect 4057 3116 4069 3122
rect 4157 3116 4169 3122
rect 4237 3116 4249 3122
rect 4298 3116 4310 3122
rect 4419 3116 4431 3122
rect 4477 3116 4489 3122
rect 4525 3116 4537 3122
rect 4587 3116 4599 3122
rect 4657 3116 4669 3122
rect 3053 2991 3060 3039
rect 3114 3033 3122 3076
rect 3220 3053 3227 3096
rect 2837 2964 2845 2970
rect 2893 2968 2923 2974
rect 2941 2964 2947 2982
rect 2827 2950 2845 2964
rect 2873 2950 2895 2962
rect 2837 2944 2845 2950
rect 2887 2944 2899 2950
rect 2941 2924 2953 2958
rect 3043 2984 3060 2991
rect 3114 2984 3122 3019
rect 3220 2991 3227 3039
rect 3320 3096 3333 3102
rect 3320 3090 3327 3096
rect 3385 3084 3392 3096
rect 3281 2992 3287 3076
rect 3371 3077 3392 3084
rect 3442 3090 3449 3096
rect 3442 3082 3453 3090
rect 3339 3066 3346 3072
rect 3407 3066 3413 3068
rect 3339 3060 3413 3066
rect 3495 3061 3503 3076
rect 3339 3052 3346 3060
rect 3300 3044 3334 3052
rect 3300 3039 3306 3044
rect 3326 3026 3353 3033
rect 3220 2984 3237 2991
rect 3143 2978 3183 2984
rect 3171 2976 3183 2978
rect 3281 2984 3343 2992
rect 3355 2988 3399 2994
rect 3337 2970 3375 2978
rect 3393 2974 3399 2988
rect 3407 2988 3413 3060
rect 3487 3047 3503 3061
rect 3473 3033 3487 3047
rect 3407 2982 3447 2988
rect 3467 2988 3481 2996
rect 3495 2984 3503 3047
rect 3337 2964 3345 2970
rect 3393 2968 3423 2974
rect 3441 2964 3447 2982
rect 3327 2950 3345 2964
rect 3373 2950 3395 2962
rect 3337 2944 3345 2950
rect 3387 2944 3399 2950
rect 3441 2924 3453 2958
rect 3560 3096 3573 3102
rect 3560 3090 3567 3096
rect 3625 3084 3632 3096
rect 3521 2992 3527 3076
rect 3611 3077 3632 3084
rect 3682 3090 3689 3096
rect 3682 3082 3693 3090
rect 3579 3066 3586 3072
rect 3647 3066 3653 3068
rect 3579 3060 3653 3066
rect 3735 3061 3743 3076
rect 3579 3052 3586 3060
rect 3540 3044 3574 3052
rect 3540 3039 3546 3044
rect 3566 3026 3593 3033
rect 3521 2984 3583 2992
rect 3595 2988 3639 2994
rect 3577 2970 3615 2978
rect 3633 2974 3639 2988
rect 3647 2988 3653 3060
rect 3727 3047 3743 3061
rect 3780 3053 3787 3096
rect 3855 3062 3863 3076
rect 3883 3076 3911 3082
rect 3871 3073 3923 3076
rect 3955 3062 3963 3076
rect 3983 3076 4011 3082
rect 3971 3073 4023 3076
rect 4049 3076 4077 3082
rect 4037 3073 4089 3076
rect 4149 3076 4177 3082
rect 4097 3062 4105 3076
rect 4137 3073 4189 3076
rect 4197 3062 4205 3076
rect 3855 3055 3880 3062
rect 3955 3055 3980 3062
rect 4080 3055 4105 3062
rect 4180 3055 4205 3062
rect 3713 3033 3727 3047
rect 3647 2982 3687 2988
rect 3707 2988 3721 2996
rect 3735 2984 3743 3047
rect 3780 2991 3787 3039
rect 3873 3033 3881 3055
rect 3973 3033 3981 3055
rect 4079 3033 4087 3055
rect 4179 3033 4187 3055
rect 4256 3041 4264 3096
rect 3780 2984 3797 2991
rect 3879 2984 3887 3019
rect 3979 2984 3987 3019
rect 4073 2984 4081 3019
rect 4173 2984 4181 3019
rect 3577 2964 3585 2970
rect 3633 2968 3663 2974
rect 3681 2964 3687 2982
rect 3567 2950 3585 2964
rect 3613 2950 3635 2962
rect 3577 2944 3585 2950
rect 3627 2944 3639 2950
rect 3681 2924 3693 2958
rect 2457 2898 2469 2904
rect 2522 2898 2534 2904
rect 2572 2898 2584 2904
rect 2639 2898 2651 2904
rect 2697 2898 2709 2904
rect 2737 2898 2749 2904
rect 2801 2898 2813 2904
rect 2867 2898 2879 2904
rect 2913 2898 2925 2904
rect 2971 2898 2983 2904
rect 3071 2898 3083 2904
rect 3151 2898 3163 2904
rect 3197 2898 3209 2904
rect 3301 2898 3313 2904
rect 3367 2898 3379 2904
rect 3413 2898 3425 2904
rect 3471 2898 3483 2904
rect 3541 2898 3553 2904
rect 3607 2898 3619 2904
rect 3653 2898 3665 2904
rect 3711 2898 3723 2904
rect 3757 2898 3769 2904
rect 3856 2898 3868 2904
rect 3906 2898 3918 2904
rect 3956 2898 3968 2904
rect 4006 2898 4018 2904
rect 4042 2898 4054 2904
rect 4092 2898 4104 2904
rect 4256 2944 4264 3027
rect 4277 3007 4283 3073
rect 4567 3096 4580 3102
rect 4451 3090 4458 3096
rect 4447 3082 4458 3090
rect 4508 3084 4515 3096
rect 4573 3090 4580 3096
rect 4397 3061 4405 3076
rect 4508 3077 4529 3084
rect 4487 3066 4493 3068
rect 4554 3066 4561 3072
rect 4346 3058 4364 3060
rect 4334 3049 4364 3058
rect 4356 3021 4364 3049
rect 4397 3047 4413 3061
rect 4487 3060 4561 3066
rect 4358 2952 4365 3007
rect 4318 2946 4365 2952
rect 4318 2944 4329 2946
rect 4142 2898 4154 2904
rect 4192 2898 4204 2904
rect 4357 2944 4365 2946
rect 4397 2984 4405 3047
rect 4413 3033 4427 3047
rect 4419 2988 4433 2996
rect 4487 2988 4493 3060
rect 4554 3052 4561 3060
rect 4566 3044 4600 3052
rect 4594 3039 4600 3044
rect 4547 3026 4574 3033
rect 4453 2982 4493 2988
rect 4501 2988 4545 2994
rect 4453 2964 4459 2982
rect 4501 2974 4507 2988
rect 4613 2992 4619 3076
rect 4649 3076 4677 3082
rect 4637 3073 4689 3076
rect 4697 3062 4705 3076
rect 4680 3055 4705 3062
rect 4679 3033 4687 3055
rect 4557 2984 4619 2992
rect 4673 2984 4681 3019
rect 4737 3007 4743 3073
rect 4477 2968 4507 2974
rect 4525 2970 4563 2978
rect 4555 2964 4563 2970
rect 4447 2924 4459 2958
rect 4505 2950 4527 2962
rect 4555 2950 4573 2964
rect 4501 2944 4513 2950
rect 4555 2944 4563 2950
rect 4237 2898 4249 2904
rect 4297 2898 4309 2904
rect 4337 2898 4349 2904
rect 4417 2898 4429 2904
rect 4475 2898 4487 2904
rect 4521 2898 4533 2904
rect 4587 2898 4599 2904
rect 4642 2898 4654 2904
rect 4692 2898 4704 2904
rect -62 2896 4776 2898
rect -62 2884 4 2896
rect -62 2882 4776 2884
rect -62 2418 -2 2882
rect 51 2876 63 2882
rect 96 2876 108 2882
rect 146 2876 158 2882
rect 197 2876 209 2882
rect 297 2876 309 2882
rect 337 2876 349 2882
rect 36 2753 44 2836
rect 189 2798 217 2804
rect 229 2870 257 2876
rect 377 2876 389 2882
rect 421 2876 433 2882
rect 496 2876 508 2882
rect 546 2876 558 2882
rect 119 2761 127 2796
rect 236 2790 248 2796
rect 221 2784 248 2790
rect 221 2761 227 2784
rect 317 2781 325 2836
rect 36 2684 44 2739
rect 113 2725 121 2747
rect 95 2718 120 2725
rect 95 2704 103 2718
rect 111 2704 163 2707
rect 213 2704 220 2747
rect 317 2718 325 2767
rect 398 2722 406 2836
rect 577 2876 589 2882
rect 617 2876 629 2882
rect 691 2876 703 2882
rect 751 2876 763 2882
rect 441 2761 449 2796
rect 519 2761 527 2796
rect 597 2781 605 2836
rect 777 2876 789 2882
rect 817 2876 829 2882
rect 857 2876 869 2882
rect 901 2876 913 2882
rect 976 2876 988 2882
rect 1026 2876 1038 2882
rect 447 2747 449 2761
rect 317 2712 341 2718
rect 329 2704 341 2712
rect 123 2698 151 2704
rect 51 2658 63 2664
rect 131 2658 143 2664
rect 180 2658 192 2664
rect 236 2658 248 2664
rect 377 2714 415 2722
rect 377 2704 389 2714
rect 441 2704 449 2747
rect 513 2725 521 2747
rect 495 2718 520 2725
rect 597 2718 605 2767
rect 676 2761 684 2796
rect 736 2761 744 2796
rect 797 2781 805 2836
rect 495 2704 503 2718
rect 597 2712 621 2718
rect 439 2694 449 2704
rect 511 2704 563 2707
rect 609 2704 621 2712
rect 676 2704 684 2747
rect 736 2704 744 2747
rect 797 2718 805 2767
rect 878 2722 886 2836
rect 1057 2876 1069 2882
rect 1097 2876 1109 2882
rect 1156 2876 1168 2882
rect 1206 2876 1218 2882
rect 1257 2876 1269 2882
rect 1315 2876 1327 2882
rect 1361 2876 1373 2882
rect 1427 2876 1439 2882
rect 1509 2876 1521 2882
rect 1581 2876 1593 2882
rect 1647 2876 1659 2882
rect 1693 2876 1705 2882
rect 1751 2876 1763 2882
rect 1802 2876 1814 2882
rect 1852 2876 1864 2882
rect 921 2761 929 2796
rect 999 2761 1007 2796
rect 1077 2781 1085 2836
rect 1287 2822 1299 2856
rect 1341 2830 1353 2836
rect 1395 2830 1403 2836
rect 1345 2818 1367 2830
rect 1395 2816 1413 2830
rect 1293 2798 1299 2816
rect 1317 2806 1347 2812
rect 1395 2810 1403 2816
rect 927 2747 929 2761
rect 797 2712 821 2718
rect 809 2704 821 2712
rect 523 2698 551 2704
rect 299 2658 311 2664
rect 407 2658 419 2664
rect 531 2658 543 2664
rect 579 2658 591 2664
rect 691 2658 703 2664
rect 751 2658 763 2664
rect 857 2714 895 2722
rect 857 2704 869 2714
rect 921 2704 929 2747
rect 993 2725 1001 2747
rect 975 2718 1000 2725
rect 1077 2718 1085 2767
rect 1179 2761 1187 2796
rect 1173 2725 1181 2747
rect 1237 2733 1245 2796
rect 1259 2784 1273 2792
rect 1293 2792 1333 2798
rect 1253 2733 1267 2747
rect 1155 2718 1180 2725
rect 1237 2719 1253 2733
rect 1327 2720 1333 2792
rect 1341 2792 1347 2806
rect 1365 2802 1403 2810
rect 1341 2786 1385 2792
rect 1397 2788 1459 2796
rect 1387 2747 1414 2754
rect 1434 2736 1440 2741
rect 1406 2728 1440 2736
rect 1394 2720 1401 2728
rect 975 2704 983 2718
rect 1077 2712 1101 2718
rect 919 2694 929 2704
rect 991 2704 1043 2707
rect 1089 2704 1101 2712
rect 1155 2704 1163 2718
rect 1003 2698 1031 2704
rect 1171 2704 1223 2707
rect 1183 2698 1211 2704
rect 1237 2704 1245 2719
rect 1327 2714 1401 2720
rect 1327 2712 1333 2714
rect 1394 2708 1401 2714
rect 1287 2690 1298 2698
rect 1291 2684 1298 2690
rect 1348 2696 1369 2703
rect 1453 2704 1459 2788
rect 1491 2761 1499 2796
rect 1535 2790 1543 2836
rect 1517 2784 1543 2790
rect 1617 2830 1625 2836
rect 1667 2830 1679 2836
rect 1607 2816 1625 2830
rect 1653 2818 1675 2830
rect 1721 2822 1733 2856
rect 1617 2810 1625 2816
rect 1617 2802 1655 2810
rect 1673 2806 1703 2812
rect 1561 2788 1623 2796
rect 1517 2778 1520 2784
rect 1491 2747 1493 2761
rect 1491 2704 1499 2747
rect 1513 2722 1520 2778
rect 1517 2716 1520 2722
rect 1517 2710 1539 2716
rect 1348 2684 1355 2696
rect 1413 2684 1420 2690
rect 1407 2678 1420 2684
rect 1531 2684 1539 2710
rect 1561 2704 1567 2788
rect 1673 2792 1679 2806
rect 1721 2798 1727 2816
rect 1635 2786 1679 2792
rect 1687 2792 1727 2798
rect 1606 2747 1633 2754
rect 1580 2736 1586 2741
rect 1580 2728 1614 2736
rect 1619 2720 1626 2728
rect 1687 2720 1693 2792
rect 1897 2876 1909 2882
rect 1957 2876 1969 2882
rect 2027 2876 2039 2882
rect 2131 2876 2143 2882
rect 2211 2876 2223 2882
rect 2291 2876 2303 2882
rect 1747 2784 1761 2792
rect 1753 2733 1767 2747
rect 1775 2733 1783 2796
rect 1833 2761 1841 2796
rect 1916 2753 1924 2836
rect 2317 2876 2329 2882
rect 2431 2876 2443 2882
rect 1619 2714 1693 2720
rect 1767 2719 1783 2733
rect 1839 2725 1847 2747
rect 1619 2708 1626 2714
rect 1687 2712 1693 2714
rect 1651 2696 1672 2703
rect 1775 2704 1783 2719
rect 1840 2718 1865 2725
rect 1600 2684 1607 2690
rect 1665 2684 1672 2696
rect 1722 2690 1733 2698
rect 1722 2684 1729 2690
rect 1600 2678 1613 2684
rect 1797 2704 1849 2707
rect 1809 2698 1837 2704
rect 1857 2704 1865 2718
rect 1916 2684 1924 2739
rect 1937 2727 1943 2773
rect 1997 2761 2005 2796
rect 2103 2789 2120 2796
rect 2183 2789 2200 2796
rect 2263 2789 2280 2796
rect 1996 2721 2004 2747
rect 2113 2741 2120 2789
rect 2193 2741 2200 2789
rect 2273 2741 2280 2789
rect 2336 2753 2344 2836
rect 2457 2876 2469 2882
rect 2517 2876 2529 2882
rect 2561 2876 2573 2882
rect 2622 2876 2634 2882
rect 2672 2876 2684 2882
rect 2403 2789 2420 2796
rect 2413 2741 2420 2789
rect 2476 2753 2484 2836
rect 1996 2714 2025 2721
rect 1957 2704 2009 2706
rect 2019 2704 2025 2714
rect 1969 2700 1997 2704
rect 2009 2664 2037 2670
rect 2113 2684 2120 2727
rect 2193 2684 2200 2727
rect 2273 2684 2280 2727
rect 2336 2684 2344 2739
rect 2413 2684 2420 2727
rect 2476 2684 2484 2739
rect 2538 2722 2546 2836
rect 2722 2876 2734 2882
rect 2772 2876 2784 2882
rect 2817 2876 2829 2882
rect 2857 2876 2869 2882
rect 2921 2876 2933 2882
rect 2987 2876 2999 2882
rect 3033 2876 3045 2882
rect 3091 2876 3103 2882
rect 3161 2876 3173 2882
rect 3227 2876 3239 2882
rect 3273 2876 3285 2882
rect 3331 2876 3343 2882
rect 3411 2876 3423 2882
rect 3491 2876 3503 2882
rect 3551 2876 3563 2882
rect 3601 2876 3613 2882
rect 3667 2876 3679 2882
rect 3713 2876 3725 2882
rect 3771 2876 3783 2882
rect 3891 2876 3903 2882
rect 3991 2876 4003 2882
rect 2581 2761 2589 2796
rect 2653 2761 2661 2796
rect 2753 2761 2761 2796
rect 2837 2781 2845 2836
rect 2957 2830 2965 2836
rect 3007 2830 3019 2836
rect 2947 2816 2965 2830
rect 2993 2818 3015 2830
rect 3061 2822 3073 2856
rect 2957 2810 2965 2816
rect 2957 2802 2995 2810
rect 3013 2806 3043 2812
rect 2901 2788 2963 2796
rect 2587 2747 2589 2761
rect 2517 2714 2555 2722
rect 2517 2704 2529 2714
rect 2581 2704 2589 2747
rect 2659 2725 2667 2747
rect 2759 2725 2767 2747
rect 2660 2718 2685 2725
rect 2760 2718 2785 2725
rect 779 2658 791 2664
rect 887 2658 899 2664
rect 1011 2658 1023 2664
rect 1059 2658 1071 2664
rect 1191 2658 1203 2664
rect 1259 2658 1271 2664
rect 1317 2658 1329 2664
rect 1365 2658 1377 2664
rect 1427 2658 1439 2664
rect 1509 2658 1521 2664
rect 1581 2658 1593 2664
rect 1643 2658 1655 2664
rect 1691 2658 1703 2664
rect 1749 2658 1761 2664
rect 1817 2658 1829 2664
rect 1897 2658 1909 2664
rect 1977 2658 1989 2664
rect 2091 2658 2103 2664
rect 2131 2658 2143 2664
rect 2171 2658 2183 2664
rect 2211 2658 2223 2664
rect 2251 2658 2263 2664
rect 2291 2658 2303 2664
rect 2317 2658 2329 2664
rect 2391 2658 2403 2664
rect 2431 2658 2443 2664
rect 2579 2694 2589 2704
rect 2617 2704 2669 2707
rect 2629 2698 2657 2704
rect 2677 2704 2685 2718
rect 2717 2704 2769 2707
rect 2729 2698 2757 2704
rect 2777 2704 2785 2718
rect 2837 2718 2845 2767
rect 2837 2712 2861 2718
rect 2849 2704 2861 2712
rect 2901 2704 2907 2788
rect 3013 2792 3019 2806
rect 3061 2798 3067 2816
rect 2975 2786 3019 2792
rect 3027 2792 3067 2798
rect 2946 2747 2973 2754
rect 2920 2736 2926 2741
rect 2920 2728 2954 2736
rect 2959 2720 2966 2728
rect 3027 2720 3033 2792
rect 3087 2784 3101 2792
rect 3093 2733 3107 2747
rect 3115 2733 3123 2796
rect 2959 2714 3033 2720
rect 3107 2719 3123 2733
rect 2959 2708 2966 2714
rect 3027 2712 3033 2714
rect 2991 2696 3012 2703
rect 3115 2704 3123 2719
rect 2940 2684 2947 2690
rect 3005 2684 3012 2696
rect 3062 2690 3073 2698
rect 3062 2684 3069 2690
rect 2940 2678 2953 2684
rect 3197 2830 3205 2836
rect 3247 2830 3259 2836
rect 3187 2816 3205 2830
rect 3233 2818 3255 2830
rect 3301 2822 3313 2856
rect 3197 2810 3205 2816
rect 3197 2802 3235 2810
rect 3253 2806 3283 2812
rect 3141 2788 3203 2796
rect 3141 2704 3147 2788
rect 3253 2792 3259 2806
rect 3301 2798 3307 2816
rect 3215 2786 3259 2792
rect 3267 2792 3307 2798
rect 3186 2747 3213 2754
rect 3160 2736 3166 2741
rect 3160 2728 3194 2736
rect 3199 2720 3206 2728
rect 3267 2720 3273 2792
rect 3327 2784 3341 2792
rect 3333 2733 3347 2747
rect 3355 2733 3363 2796
rect 3396 2753 3404 2836
rect 3637 2830 3645 2836
rect 3687 2830 3699 2836
rect 3627 2816 3645 2830
rect 3673 2818 3695 2830
rect 3741 2822 3753 2856
rect 3637 2810 3645 2816
rect 3637 2802 3675 2810
rect 3693 2806 3723 2812
rect 3463 2789 3480 2796
rect 3473 2741 3480 2789
rect 3536 2761 3544 2796
rect 3581 2788 3643 2796
rect 3199 2714 3273 2720
rect 3347 2719 3363 2733
rect 3199 2708 3206 2714
rect 3267 2712 3273 2714
rect 3231 2696 3252 2703
rect 3355 2704 3363 2719
rect 3180 2684 3187 2690
rect 3245 2684 3252 2696
rect 3302 2690 3313 2698
rect 3302 2684 3309 2690
rect 3180 2678 3193 2684
rect 3396 2684 3404 2739
rect 3473 2684 3480 2727
rect 3536 2704 3544 2747
rect 3581 2704 3587 2788
rect 3693 2792 3699 2806
rect 3741 2798 3747 2816
rect 3655 2786 3699 2792
rect 3707 2792 3747 2798
rect 3626 2747 3653 2754
rect 3600 2736 3606 2741
rect 3600 2728 3634 2736
rect 3639 2720 3646 2728
rect 3707 2720 3713 2792
rect 3843 2870 3871 2876
rect 3883 2798 3911 2804
rect 4022 2876 4034 2882
rect 4072 2876 4084 2882
rect 4136 2876 4148 2882
rect 4186 2876 4198 2882
rect 4217 2876 4229 2882
rect 4321 2876 4333 2882
rect 4387 2876 4399 2882
rect 4433 2876 4445 2882
rect 4491 2876 4503 2882
rect 4542 2876 4554 2882
rect 4592 2876 4604 2882
rect 3767 2784 3781 2792
rect 3773 2733 3787 2747
rect 3795 2733 3803 2796
rect 3852 2790 3864 2796
rect 3852 2784 3879 2790
rect 3963 2789 3980 2796
rect 3873 2761 3879 2784
rect 3639 2714 3713 2720
rect 3787 2719 3803 2733
rect 3639 2708 3646 2714
rect 3707 2712 3713 2714
rect 2457 2658 2469 2664
rect 2547 2658 2559 2664
rect 2637 2658 2649 2664
rect 2737 2658 2749 2664
rect 2819 2658 2831 2664
rect 2921 2658 2933 2664
rect 2983 2658 2995 2664
rect 3031 2658 3043 2664
rect 3089 2658 3101 2664
rect 3161 2658 3173 2664
rect 3223 2658 3235 2664
rect 3271 2658 3283 2664
rect 3329 2658 3341 2664
rect 3411 2658 3423 2664
rect 3671 2696 3692 2703
rect 3795 2704 3803 2719
rect 3880 2704 3887 2747
rect 3973 2741 3980 2789
rect 4053 2761 4061 2796
rect 4159 2761 4167 2796
rect 4240 2789 4257 2796
rect 4357 2830 4365 2836
rect 4407 2830 4419 2836
rect 4347 2816 4365 2830
rect 4393 2818 4415 2830
rect 4461 2822 4473 2856
rect 4357 2810 4365 2816
rect 4357 2802 4395 2810
rect 4413 2806 4443 2812
rect 3620 2684 3627 2690
rect 3685 2684 3692 2696
rect 3742 2690 3753 2698
rect 3742 2684 3749 2690
rect 3620 2678 3633 2684
rect 3973 2684 3980 2727
rect 4059 2725 4067 2747
rect 4153 2725 4161 2747
rect 4240 2741 4247 2789
rect 4301 2788 4363 2796
rect 4060 2718 4085 2725
rect 4017 2704 4069 2707
rect 3451 2658 3463 2664
rect 3491 2658 3503 2664
rect 3551 2658 3563 2664
rect 3601 2658 3613 2664
rect 3663 2658 3675 2664
rect 3711 2658 3723 2664
rect 3769 2658 3781 2664
rect 3852 2658 3864 2664
rect 3908 2658 3920 2664
rect 4029 2698 4057 2704
rect 4077 2704 4085 2718
rect 4135 2718 4160 2725
rect 4135 2704 4143 2718
rect 4151 2704 4203 2707
rect 4163 2698 4191 2704
rect 4240 2684 4247 2727
rect 4301 2704 4307 2788
rect 4413 2792 4419 2806
rect 4461 2798 4467 2816
rect 4375 2786 4419 2792
rect 4427 2792 4467 2798
rect 4346 2747 4373 2754
rect 4320 2736 4326 2741
rect 4320 2728 4354 2736
rect 4359 2720 4366 2728
rect 4427 2720 4433 2792
rect 4637 2876 4649 2882
rect 4677 2876 4689 2882
rect 4487 2784 4501 2792
rect 4493 2733 4507 2747
rect 4515 2733 4523 2796
rect 4573 2761 4581 2796
rect 4657 2781 4665 2836
rect 4359 2714 4433 2720
rect 4507 2719 4523 2733
rect 4579 2725 4587 2747
rect 4359 2708 4366 2714
rect 4427 2712 4433 2714
rect 4391 2696 4412 2703
rect 4515 2704 4523 2719
rect 4580 2718 4605 2725
rect 4340 2684 4347 2690
rect 4405 2684 4412 2696
rect 4462 2690 4473 2698
rect 4462 2684 4469 2690
rect 4340 2678 4353 2684
rect 4537 2704 4589 2707
rect 4549 2698 4577 2704
rect 4597 2704 4605 2718
rect 4657 2718 4665 2767
rect 4657 2712 4681 2718
rect 4669 2704 4681 2712
rect 3951 2658 3963 2664
rect 3991 2658 4003 2664
rect 4037 2658 4049 2664
rect 4171 2658 4183 2664
rect 4217 2658 4229 2664
rect 4257 2658 4269 2664
rect 4321 2658 4333 2664
rect 4383 2658 4395 2664
rect 4431 2658 4443 2664
rect 4489 2658 4501 2664
rect 4557 2658 4569 2664
rect 4639 2658 4651 2664
rect 4782 2658 4842 3122
rect 4 2656 4842 2658
rect 4776 2644 4842 2656
rect 4 2642 4842 2644
rect 18 2636 30 2642
rect 120 2636 132 2642
rect 170 2636 182 2642
rect 251 2636 263 2642
rect 321 2636 333 2642
rect 398 2636 410 2642
rect 448 2636 460 2642
rect 550 2636 562 2642
rect 631 2636 643 2642
rect 711 2636 723 2642
rect 789 2636 801 2642
rect 890 2636 902 2642
rect 971 2636 983 2642
rect 1019 2636 1031 2642
rect 1170 2636 1182 2642
rect 1231 2636 1243 2642
rect 1311 2636 1323 2642
rect 1359 2636 1371 2642
rect 1437 2636 1449 2642
rect 1549 2636 1561 2642
rect 1601 2636 1613 2642
rect 1663 2636 1675 2642
rect 1711 2636 1723 2642
rect 1769 2636 1781 2642
rect 1819 2636 1831 2642
rect 1899 2636 1911 2642
rect 1978 2636 1990 2642
rect 2077 2636 2089 2642
rect 2117 2636 2129 2642
rect 2191 2636 2203 2642
rect 160 2596 186 2607
rect 66 2578 84 2580
rect 54 2569 84 2578
rect 76 2541 84 2569
rect 178 2553 186 2596
rect 236 2561 244 2616
rect 291 2596 301 2606
rect 291 2553 299 2596
rect 351 2586 363 2596
rect 325 2578 363 2586
rect 394 2596 420 2607
rect 477 2597 493 2603
rect 78 2472 85 2527
rect 178 2504 186 2539
rect 38 2466 85 2472
rect 38 2464 49 2466
rect 77 2464 85 2466
rect 117 2498 157 2504
rect 117 2496 129 2498
rect 236 2464 244 2547
rect 291 2539 293 2553
rect 291 2504 299 2539
rect 334 2464 342 2578
rect 394 2553 402 2596
rect 394 2504 402 2539
rect 477 2523 483 2597
rect 496 2578 514 2580
rect 496 2569 526 2578
rect 595 2582 603 2596
rect 623 2596 651 2602
rect 611 2593 663 2596
rect 595 2575 620 2582
rect 496 2541 504 2569
rect 547 2557 593 2563
rect 613 2553 621 2575
rect 696 2553 704 2596
rect 759 2588 771 2596
rect 759 2582 783 2588
rect 467 2517 483 2523
rect 423 2498 463 2504
rect 451 2496 463 2498
rect 495 2472 502 2527
rect 619 2504 627 2539
rect 696 2504 704 2539
rect 775 2533 783 2582
rect 807 2577 823 2583
rect 495 2466 542 2472
rect 495 2464 503 2466
rect 531 2464 542 2466
rect 17 2418 29 2424
rect 57 2418 69 2424
rect 137 2418 149 2424
rect 251 2418 263 2424
rect 307 2418 319 2424
rect 351 2418 363 2424
rect 431 2418 443 2424
rect 511 2418 523 2424
rect 551 2418 563 2424
rect 775 2464 783 2519
rect 817 2503 823 2577
rect 836 2578 854 2580
rect 836 2569 866 2578
rect 935 2582 943 2596
rect 963 2596 991 2602
rect 951 2593 1003 2596
rect 1049 2588 1061 2596
rect 1037 2582 1061 2588
rect 935 2575 960 2582
rect 836 2541 844 2569
rect 953 2553 961 2575
rect 807 2497 823 2503
rect 835 2472 842 2527
rect 959 2504 967 2539
rect 1037 2533 1045 2582
rect 1116 2578 1134 2580
rect 1116 2569 1146 2578
rect 1116 2541 1124 2569
rect 1216 2561 1224 2616
rect 1275 2582 1283 2596
rect 1303 2596 1331 2602
rect 1620 2616 1633 2622
rect 1620 2610 1627 2616
rect 1685 2604 1692 2616
rect 1291 2593 1343 2596
rect 1389 2588 1401 2596
rect 1377 2582 1401 2588
rect 1275 2575 1300 2582
rect 1293 2553 1301 2575
rect 835 2466 882 2472
rect 835 2464 843 2466
rect 596 2418 608 2424
rect 646 2418 658 2424
rect 711 2418 723 2424
rect 871 2464 882 2466
rect 751 2418 763 2424
rect 791 2418 803 2424
rect 851 2418 863 2424
rect 891 2418 903 2424
rect 1037 2464 1045 2519
rect 1115 2472 1122 2527
rect 1115 2466 1162 2472
rect 1115 2464 1123 2466
rect 936 2418 948 2424
rect 986 2418 998 2424
rect 1151 2464 1162 2466
rect 1216 2464 1224 2547
rect 1299 2504 1307 2539
rect 1377 2533 1385 2582
rect 1456 2553 1464 2596
rect 1519 2588 1531 2596
rect 1519 2582 1543 2588
rect 1017 2418 1029 2424
rect 1057 2418 1069 2424
rect 1131 2418 1143 2424
rect 1171 2418 1183 2424
rect 1231 2418 1243 2424
rect 1377 2464 1385 2519
rect 1456 2504 1464 2539
rect 1535 2533 1543 2582
rect 1276 2418 1288 2424
rect 1326 2418 1338 2424
rect 1357 2418 1369 2424
rect 1397 2418 1409 2424
rect 1535 2464 1543 2519
rect 1581 2512 1587 2596
rect 1671 2597 1692 2604
rect 1742 2610 1749 2616
rect 1742 2602 1753 2610
rect 1639 2586 1646 2592
rect 1707 2586 1713 2588
rect 1639 2580 1713 2586
rect 1795 2581 1803 2596
rect 1849 2588 1861 2596
rect 1929 2588 1941 2596
rect 1639 2572 1646 2580
rect 1600 2564 1634 2572
rect 1600 2559 1606 2564
rect 1626 2546 1653 2553
rect 1581 2504 1643 2512
rect 1655 2508 1699 2514
rect 1637 2490 1675 2498
rect 1693 2494 1699 2508
rect 1707 2508 1713 2580
rect 1787 2567 1803 2581
rect 1773 2553 1787 2567
rect 1707 2502 1747 2508
rect 1767 2508 1781 2516
rect 1795 2504 1803 2567
rect 1837 2582 1861 2588
rect 1917 2582 1941 2588
rect 1837 2533 1845 2582
rect 1917 2533 1925 2582
rect 2231 2636 2243 2642
rect 2271 2636 2283 2642
rect 2331 2636 2343 2642
rect 2411 2636 2423 2642
rect 2457 2636 2469 2642
rect 2497 2636 2509 2642
rect 2567 2636 2579 2642
rect 2657 2636 2669 2642
rect 2789 2636 2801 2642
rect 2026 2578 2044 2580
rect 2014 2569 2044 2578
rect 2100 2573 2107 2616
rect 2036 2541 2044 2569
rect 2176 2561 2184 2616
rect 2253 2573 2260 2616
rect 1637 2484 1645 2490
rect 1693 2488 1723 2494
rect 1741 2484 1747 2502
rect 1627 2470 1645 2484
rect 1673 2470 1695 2482
rect 1637 2464 1645 2470
rect 1687 2464 1699 2470
rect 1741 2444 1753 2478
rect 1837 2464 1845 2519
rect 1917 2464 1925 2519
rect 2038 2472 2045 2527
rect 2100 2511 2107 2559
rect 2316 2561 2324 2616
rect 2375 2582 2383 2596
rect 2403 2596 2431 2602
rect 2391 2593 2443 2596
rect 2375 2575 2400 2582
rect 2100 2504 2117 2511
rect 1998 2466 2045 2472
rect 1998 2464 2009 2466
rect 1437 2418 1449 2424
rect 1511 2418 1523 2424
rect 1551 2418 1563 2424
rect 1601 2418 1613 2424
rect 1667 2418 1679 2424
rect 1713 2418 1725 2424
rect 1771 2418 1783 2424
rect 1817 2418 1829 2424
rect 1857 2418 1869 2424
rect 1897 2418 1909 2424
rect 1937 2418 1949 2424
rect 2037 2464 2045 2466
rect 2176 2464 2184 2547
rect 2253 2511 2260 2559
rect 2393 2553 2401 2575
rect 2480 2573 2487 2616
rect 2599 2596 2609 2606
rect 2537 2586 2549 2596
rect 2537 2578 2575 2586
rect 2243 2504 2260 2511
rect 2316 2464 2324 2547
rect 2399 2504 2407 2539
rect 2480 2511 2487 2559
rect 2480 2504 2497 2511
rect 1977 2418 1989 2424
rect 2017 2418 2029 2424
rect 2077 2418 2089 2424
rect 2191 2418 2203 2424
rect 2271 2418 2283 2424
rect 2331 2418 2343 2424
rect 2376 2418 2388 2424
rect 2426 2418 2438 2424
rect 2558 2464 2566 2578
rect 2601 2553 2609 2596
rect 2649 2596 2677 2602
rect 2637 2593 2689 2596
rect 2817 2636 2825 2642
rect 2857 2636 2869 2642
rect 2919 2636 2931 2642
rect 3019 2636 3031 2642
rect 3097 2636 3109 2642
rect 3209 2636 3221 2642
rect 3309 2636 3321 2642
rect 2697 2582 2705 2596
rect 2759 2588 2771 2596
rect 2843 2588 2849 2616
rect 2759 2582 2783 2588
rect 2843 2582 2853 2588
rect 2680 2575 2705 2582
rect 2607 2539 2609 2553
rect 2679 2553 2687 2575
rect 2601 2504 2609 2539
rect 2673 2504 2681 2539
rect 2775 2533 2783 2582
rect 2858 2521 2864 2576
rect 2880 2561 2887 2596
rect 2949 2588 2961 2596
rect 2937 2582 2961 2588
rect 3001 2590 3009 2616
rect 3089 2596 3117 2602
rect 3001 2584 3023 2590
rect 2775 2464 2783 2519
rect 2817 2512 2853 2520
rect 2817 2504 2825 2512
rect 2457 2418 2469 2424
rect 2537 2418 2549 2424
rect 2581 2418 2593 2424
rect 2642 2418 2654 2424
rect 2692 2418 2704 2424
rect 2874 2503 2883 2547
rect 2937 2533 2945 2582
rect 3020 2578 3023 2584
rect 3020 2522 3027 2578
rect 3041 2553 3049 2596
rect 3077 2593 3129 2596
rect 3137 2582 3145 2596
rect 3120 2575 3145 2582
rect 3047 2539 3049 2553
rect 3119 2553 3127 2575
rect 3191 2553 3199 2596
rect 3231 2590 3239 2616
rect 3217 2584 3239 2590
rect 3340 2636 3352 2642
rect 3396 2636 3408 2642
rect 3479 2636 3491 2642
rect 3569 2636 3581 2642
rect 3641 2636 3653 2642
rect 3703 2636 3715 2642
rect 3751 2636 3763 2642
rect 3809 2636 3821 2642
rect 3878 2636 3890 2642
rect 3928 2636 3940 2642
rect 3279 2588 3291 2596
rect 3217 2578 3220 2584
rect 3279 2582 3303 2588
rect 3191 2539 3193 2553
rect 2879 2494 2883 2503
rect 2937 2464 2945 2519
rect 3020 2516 3023 2522
rect 2997 2510 3023 2516
rect 2997 2464 3005 2510
rect 3041 2504 3049 2539
rect 3113 2504 3121 2539
rect 3191 2504 3199 2539
rect 3213 2522 3220 2578
rect 3295 2533 3303 2582
rect 3217 2516 3220 2522
rect 3373 2553 3380 2596
rect 3461 2590 3469 2616
rect 3461 2584 3483 2590
rect 3480 2578 3483 2584
rect 3217 2510 3243 2516
rect 3235 2464 3243 2510
rect 3295 2464 3303 2519
rect 3381 2516 3387 2539
rect 3480 2522 3487 2578
rect 3501 2553 3509 2596
rect 3507 2539 3509 2553
rect 3480 2516 3483 2522
rect 3381 2510 3408 2516
rect 3396 2504 3408 2510
rect 3457 2510 3483 2516
rect 3349 2496 3377 2502
rect 3389 2424 3417 2430
rect 3457 2464 3465 2510
rect 3501 2504 3509 2539
rect 3551 2553 3559 2596
rect 3591 2590 3599 2616
rect 3577 2584 3599 2590
rect 3660 2616 3673 2622
rect 3660 2610 3667 2616
rect 3725 2604 3732 2616
rect 3577 2578 3580 2584
rect 3551 2539 3553 2553
rect 3551 2504 3559 2539
rect 3573 2522 3580 2578
rect 3577 2516 3580 2522
rect 3577 2510 3603 2516
rect 3595 2464 3603 2510
rect 3621 2512 3627 2596
rect 3711 2597 3732 2604
rect 3782 2610 3789 2616
rect 3782 2602 3793 2610
rect 3679 2586 3686 2592
rect 3747 2586 3753 2588
rect 3679 2580 3753 2586
rect 3835 2581 3843 2596
rect 3679 2572 3686 2580
rect 3640 2564 3674 2572
rect 3640 2559 3646 2564
rect 3666 2546 3693 2553
rect 3621 2504 3683 2512
rect 3695 2508 3739 2514
rect 3677 2490 3715 2498
rect 3733 2494 3739 2508
rect 3747 2508 3753 2580
rect 3827 2567 3843 2581
rect 3813 2553 3827 2567
rect 3747 2502 3787 2508
rect 3807 2508 3821 2516
rect 3835 2504 3843 2567
rect 3874 2596 3900 2607
rect 3957 2636 3969 2642
rect 3997 2636 4009 2642
rect 4037 2636 4049 2642
rect 4077 2636 4089 2642
rect 4117 2636 4129 2642
rect 4157 2636 4169 2642
rect 4197 2636 4209 2642
rect 4261 2636 4273 2642
rect 4323 2636 4335 2642
rect 4371 2636 4383 2642
rect 4429 2636 4441 2642
rect 4497 2636 4509 2642
rect 4579 2636 4591 2642
rect 4659 2636 4671 2642
rect 3874 2553 3882 2596
rect 3980 2573 3987 2616
rect 4280 2616 4293 2622
rect 4280 2610 4287 2616
rect 4345 2604 4352 2616
rect 4056 2590 4068 2596
rect 4097 2590 4109 2596
rect 4136 2590 4148 2596
rect 4176 2590 4188 2596
rect 4056 2582 4083 2590
rect 4097 2582 4122 2590
rect 4136 2582 4162 2590
rect 4176 2589 4194 2590
rect 4176 2582 4195 2589
rect 4075 2576 4083 2582
rect 4114 2576 4122 2582
rect 4154 2576 4162 2582
rect 4075 2564 4090 2576
rect 4114 2564 4130 2576
rect 4154 2564 4170 2576
rect 3874 2504 3882 2539
rect 3980 2511 3987 2559
rect 4075 2518 4083 2564
rect 4114 2518 4122 2564
rect 4154 2518 4162 2564
rect 4188 2561 4195 2582
rect 4188 2547 4193 2561
rect 4188 2518 4195 2547
rect 3980 2504 3997 2511
rect 4057 2510 4083 2518
rect 4097 2510 4122 2518
rect 4137 2510 4162 2518
rect 4177 2510 4195 2518
rect 4241 2512 4247 2596
rect 4331 2597 4352 2604
rect 4402 2610 4409 2616
rect 4402 2602 4413 2610
rect 4299 2586 4306 2592
rect 4367 2586 4373 2588
rect 4299 2580 4373 2586
rect 4455 2581 4463 2596
rect 4489 2596 4517 2602
rect 4477 2593 4529 2596
rect 4537 2582 4545 2596
rect 4609 2588 4621 2596
rect 4689 2588 4701 2596
rect 4299 2572 4306 2580
rect 4260 2564 4294 2572
rect 4260 2559 4266 2564
rect 4286 2546 4313 2553
rect 4057 2504 4069 2510
rect 4097 2504 4109 2510
rect 4137 2504 4149 2510
rect 4177 2504 4189 2510
rect 4241 2504 4303 2512
rect 4315 2508 4359 2514
rect 3677 2484 3685 2490
rect 3733 2488 3763 2494
rect 3781 2484 3787 2502
rect 3667 2470 3685 2484
rect 3713 2470 3735 2482
rect 3677 2464 3685 2470
rect 3727 2464 3739 2470
rect 3781 2444 3793 2478
rect 3903 2498 3943 2504
rect 3931 2496 3943 2498
rect 4297 2490 4335 2498
rect 4353 2494 4359 2508
rect 4367 2508 4373 2580
rect 4447 2567 4463 2581
rect 4520 2575 4545 2582
rect 4597 2582 4621 2588
rect 4677 2582 4701 2588
rect 4433 2553 4447 2567
rect 4367 2502 4407 2508
rect 4427 2508 4441 2516
rect 4455 2504 4463 2567
rect 4519 2553 4527 2575
rect 4513 2504 4521 2539
rect 4597 2533 4605 2582
rect 4677 2533 4685 2582
rect 4297 2484 4305 2490
rect 4353 2488 4383 2494
rect 4401 2484 4407 2502
rect 4287 2470 4305 2484
rect 4333 2470 4355 2482
rect 4297 2464 4305 2470
rect 4347 2464 4359 2470
rect 4401 2444 4413 2478
rect 4597 2464 4605 2519
rect 4677 2464 4685 2519
rect 2751 2418 2763 2424
rect 2791 2418 2803 2424
rect 2847 2418 2859 2424
rect 2917 2418 2929 2424
rect 2957 2418 2969 2424
rect 3019 2418 3031 2424
rect 3082 2418 3094 2424
rect 3132 2418 3144 2424
rect 3209 2418 3221 2424
rect 3271 2418 3283 2424
rect 3311 2418 3323 2424
rect 3357 2418 3369 2424
rect 3479 2418 3491 2424
rect 3569 2418 3581 2424
rect 3641 2418 3653 2424
rect 3707 2418 3719 2424
rect 3753 2418 3765 2424
rect 3811 2418 3823 2424
rect 3911 2418 3923 2424
rect 3957 2418 3969 2424
rect 4037 2418 4049 2424
rect 4077 2418 4089 2424
rect 4117 2418 4129 2424
rect 4157 2418 4169 2424
rect 4197 2418 4209 2424
rect 4261 2418 4273 2424
rect 4327 2418 4339 2424
rect 4373 2418 4385 2424
rect 4431 2418 4443 2424
rect 4482 2418 4494 2424
rect 4532 2418 4544 2424
rect 4577 2418 4589 2424
rect 4617 2418 4629 2424
rect 4657 2418 4669 2424
rect 4697 2418 4709 2424
rect -62 2416 4776 2418
rect -62 2404 4 2416
rect -62 2402 4776 2404
rect -62 1938 -2 2402
rect 51 2396 63 2402
rect 91 2396 103 2402
rect 35 2354 43 2356
rect 136 2396 148 2402
rect 186 2396 198 2402
rect 71 2354 82 2356
rect 35 2348 82 2354
rect 35 2293 42 2348
rect 117 2337 133 2343
rect 36 2251 44 2279
rect 117 2263 123 2337
rect 222 2396 234 2402
rect 272 2396 284 2402
rect 317 2396 329 2402
rect 357 2396 369 2402
rect 437 2396 449 2402
rect 522 2396 534 2402
rect 572 2396 584 2402
rect 671 2396 683 2402
rect 717 2396 729 2402
rect 807 2396 819 2402
rect 851 2396 863 2402
rect 338 2354 349 2356
rect 377 2354 385 2356
rect 338 2348 385 2354
rect 159 2281 167 2316
rect 253 2281 261 2316
rect 378 2293 385 2348
rect 417 2322 429 2324
rect 417 2316 457 2322
rect 691 2322 703 2324
rect 663 2316 703 2322
rect 107 2257 123 2263
rect 36 2242 66 2251
rect 153 2245 161 2267
rect 478 2281 486 2316
rect 553 2281 561 2316
rect 634 2281 642 2316
rect 259 2245 267 2267
rect 376 2251 384 2279
rect 36 2240 54 2242
rect 135 2238 160 2245
rect 260 2238 285 2245
rect 135 2224 143 2238
rect 151 2224 203 2227
rect 163 2218 191 2224
rect 217 2224 269 2227
rect 229 2218 257 2224
rect 277 2224 285 2238
rect 354 2242 384 2251
rect 366 2240 384 2242
rect 478 2224 486 2267
rect 736 2273 744 2356
rect 877 2396 889 2402
rect 917 2396 929 2402
rect 957 2396 969 2402
rect 1001 2396 1013 2402
rect 1076 2396 1088 2402
rect 1126 2396 1138 2402
rect 791 2281 799 2316
rect 559 2245 567 2267
rect 560 2238 585 2245
rect 460 2213 486 2224
rect 517 2224 569 2227
rect 529 2218 557 2224
rect 577 2224 585 2238
rect 634 2224 642 2267
rect 791 2267 793 2281
rect 634 2213 660 2224
rect 736 2204 744 2259
rect 791 2224 799 2267
rect 834 2242 842 2356
rect 897 2301 905 2356
rect 825 2234 863 2242
rect 851 2224 863 2234
rect 897 2238 905 2287
rect 978 2242 986 2356
rect 1176 2396 1188 2402
rect 1226 2396 1238 2402
rect 1281 2396 1293 2402
rect 1347 2396 1359 2402
rect 1393 2396 1405 2402
rect 1451 2396 1463 2402
rect 1516 2396 1528 2402
rect 1566 2396 1578 2402
rect 1621 2396 1633 2402
rect 1687 2396 1699 2402
rect 1733 2396 1745 2402
rect 1791 2396 1803 2402
rect 1871 2396 1883 2402
rect 1931 2396 1943 2402
rect 1317 2350 1325 2356
rect 1367 2350 1379 2356
rect 1307 2336 1325 2350
rect 1353 2338 1375 2350
rect 1421 2342 1433 2376
rect 1317 2330 1325 2336
rect 1317 2322 1355 2330
rect 1373 2326 1403 2332
rect 1021 2281 1029 2316
rect 1099 2281 1107 2316
rect 1199 2281 1207 2316
rect 1261 2308 1323 2316
rect 1027 2267 1029 2281
rect 897 2232 921 2238
rect 909 2224 921 2232
rect 791 2214 801 2224
rect 90 2178 102 2184
rect 171 2178 183 2184
rect 237 2178 249 2184
rect 318 2178 330 2184
rect 420 2178 432 2184
rect 470 2178 482 2184
rect 537 2178 549 2184
rect 638 2178 650 2184
rect 688 2178 700 2184
rect 957 2234 995 2242
rect 957 2224 969 2234
rect 1021 2224 1029 2267
rect 1093 2245 1101 2267
rect 1193 2245 1201 2267
rect 1075 2238 1100 2245
rect 1175 2238 1200 2245
rect 1075 2224 1083 2238
rect 1019 2214 1029 2224
rect 1091 2224 1143 2227
rect 1175 2224 1183 2238
rect 1103 2218 1131 2224
rect 1191 2224 1243 2227
rect 1203 2218 1231 2224
rect 1261 2224 1267 2308
rect 1373 2312 1379 2326
rect 1421 2318 1427 2336
rect 1335 2306 1379 2312
rect 1387 2312 1427 2318
rect 1306 2267 1333 2274
rect 1280 2256 1286 2261
rect 1280 2248 1314 2256
rect 1319 2240 1326 2248
rect 1387 2240 1393 2312
rect 1657 2350 1665 2356
rect 1707 2350 1719 2356
rect 1647 2336 1665 2350
rect 1693 2338 1715 2350
rect 1761 2342 1773 2376
rect 1657 2330 1665 2336
rect 1657 2322 1695 2330
rect 1713 2326 1743 2332
rect 1447 2304 1461 2312
rect 1453 2253 1467 2267
rect 1475 2253 1483 2316
rect 1539 2281 1547 2316
rect 1601 2308 1663 2316
rect 1319 2234 1393 2240
rect 1467 2239 1483 2253
rect 1533 2245 1541 2267
rect 1319 2228 1326 2234
rect 1387 2232 1393 2234
rect 1351 2216 1372 2223
rect 1475 2224 1483 2239
rect 1515 2238 1540 2245
rect 1515 2224 1523 2238
rect 1300 2204 1307 2210
rect 1365 2204 1372 2216
rect 1422 2210 1433 2218
rect 1422 2204 1429 2210
rect 1300 2198 1313 2204
rect 1531 2224 1583 2227
rect 1543 2218 1571 2224
rect 1601 2224 1607 2308
rect 1713 2312 1719 2326
rect 1761 2318 1767 2336
rect 1675 2306 1719 2312
rect 1727 2312 1767 2318
rect 1646 2267 1673 2274
rect 1620 2256 1626 2261
rect 1620 2248 1654 2256
rect 1659 2240 1666 2248
rect 1727 2240 1733 2312
rect 1962 2396 1974 2402
rect 2012 2396 2024 2402
rect 2081 2396 2093 2402
rect 2147 2396 2159 2402
rect 2193 2396 2205 2402
rect 2251 2396 2263 2402
rect 2351 2396 2363 2402
rect 2451 2396 2463 2402
rect 2497 2396 2509 2402
rect 2537 2396 2549 2402
rect 2597 2396 2609 2402
rect 2641 2396 2653 2402
rect 2717 2396 2729 2402
rect 2775 2396 2787 2402
rect 2821 2396 2833 2402
rect 2887 2396 2899 2402
rect 2956 2396 2968 2402
rect 3006 2396 3018 2402
rect 1787 2304 1801 2312
rect 1793 2253 1807 2267
rect 1815 2253 1823 2316
rect 1856 2273 1864 2356
rect 1916 2273 1924 2356
rect 2117 2350 2125 2356
rect 2167 2350 2179 2356
rect 2107 2336 2125 2350
rect 2153 2338 2175 2350
rect 2221 2342 2233 2376
rect 2117 2330 2125 2336
rect 2117 2322 2155 2330
rect 2173 2326 2203 2332
rect 1993 2281 2001 2316
rect 2061 2308 2123 2316
rect 1659 2234 1733 2240
rect 1807 2239 1823 2253
rect 1659 2228 1666 2234
rect 1727 2232 1733 2234
rect 1691 2216 1712 2223
rect 1815 2224 1823 2239
rect 1640 2204 1647 2210
rect 1705 2204 1712 2216
rect 1762 2210 1773 2218
rect 1762 2204 1769 2210
rect 1640 2198 1653 2204
rect 1856 2204 1864 2259
rect 1916 2204 1924 2259
rect 1999 2245 2007 2267
rect 2000 2238 2025 2245
rect 1957 2224 2009 2227
rect 1969 2218 1997 2224
rect 2017 2224 2025 2238
rect 2061 2224 2067 2308
rect 2173 2312 2179 2326
rect 2221 2318 2227 2336
rect 2135 2306 2179 2312
rect 2187 2312 2227 2318
rect 2106 2267 2133 2274
rect 2080 2256 2086 2261
rect 2080 2248 2114 2256
rect 2119 2240 2126 2248
rect 2187 2240 2193 2312
rect 2371 2322 2383 2324
rect 2343 2316 2383 2322
rect 2518 2354 2529 2356
rect 2557 2354 2565 2356
rect 2518 2348 2565 2354
rect 2471 2322 2483 2324
rect 2443 2316 2483 2322
rect 2247 2304 2261 2312
rect 2253 2253 2267 2267
rect 2275 2253 2283 2316
rect 2314 2281 2322 2316
rect 2414 2281 2422 2316
rect 2558 2293 2565 2348
rect 2119 2234 2193 2240
rect 2267 2239 2283 2253
rect 2119 2228 2126 2234
rect 2187 2232 2193 2234
rect 2151 2216 2172 2223
rect 2275 2224 2283 2239
rect 2100 2204 2107 2210
rect 2165 2204 2172 2216
rect 2222 2210 2233 2218
rect 2222 2204 2229 2210
rect 2100 2198 2113 2204
rect 2314 2224 2322 2267
rect 2414 2224 2422 2267
rect 2556 2251 2564 2279
rect 2314 2213 2340 2224
rect 2414 2213 2440 2224
rect 717 2178 729 2184
rect 821 2178 833 2184
rect 879 2178 891 2184
rect 987 2178 999 2184
rect 1111 2178 1123 2184
rect 1211 2178 1223 2184
rect 1281 2178 1293 2184
rect 1343 2178 1355 2184
rect 1391 2178 1403 2184
rect 1449 2178 1461 2184
rect 1551 2178 1563 2184
rect 1621 2178 1633 2184
rect 1683 2178 1695 2184
rect 1731 2178 1743 2184
rect 1789 2178 1801 2184
rect 1871 2178 1883 2184
rect 1931 2178 1943 2184
rect 1977 2178 1989 2184
rect 2081 2178 2093 2184
rect 2143 2178 2155 2184
rect 2191 2178 2203 2184
rect 2249 2178 2261 2184
rect 2318 2178 2330 2184
rect 2368 2178 2380 2184
rect 2418 2178 2430 2184
rect 2468 2178 2480 2184
rect 2534 2242 2564 2251
rect 2618 2242 2626 2356
rect 2747 2342 2759 2376
rect 2801 2350 2813 2356
rect 2855 2350 2863 2356
rect 2805 2338 2827 2350
rect 2855 2336 2873 2350
rect 2753 2318 2759 2336
rect 2777 2326 2807 2332
rect 2855 2330 2863 2336
rect 2661 2281 2669 2316
rect 2667 2267 2669 2281
rect 2546 2240 2564 2242
rect 2597 2234 2635 2242
rect 2597 2224 2609 2234
rect 2661 2224 2669 2267
rect 2659 2214 2669 2224
rect 2697 2253 2705 2316
rect 2719 2304 2733 2312
rect 2753 2312 2793 2318
rect 2713 2253 2727 2267
rect 2697 2239 2713 2253
rect 2787 2240 2793 2312
rect 2801 2312 2807 2326
rect 2825 2322 2863 2330
rect 3056 2396 3068 2402
rect 3106 2396 3118 2402
rect 3142 2396 3154 2402
rect 3192 2396 3204 2402
rect 3257 2396 3269 2402
rect 3315 2396 3327 2402
rect 3361 2396 3373 2402
rect 3427 2396 3439 2402
rect 3496 2396 3508 2402
rect 3546 2396 3558 2402
rect 3631 2396 3643 2402
rect 3687 2396 3699 2402
rect 3771 2396 3783 2402
rect 3811 2396 3823 2402
rect 3911 2396 3923 2402
rect 4031 2396 4043 2402
rect 4101 2396 4113 2402
rect 4167 2396 4179 2402
rect 4213 2396 4225 2402
rect 4271 2396 4283 2402
rect 4337 2396 4349 2402
rect 4395 2396 4407 2402
rect 4441 2396 4453 2402
rect 4507 2396 4519 2402
rect 4562 2396 4574 2402
rect 4612 2396 4624 2402
rect 3287 2342 3299 2376
rect 3341 2350 3353 2356
rect 3395 2350 3403 2356
rect 3345 2338 3367 2350
rect 3395 2336 3413 2350
rect 3293 2318 3299 2336
rect 3317 2326 3347 2332
rect 3395 2330 3403 2336
rect 2801 2306 2845 2312
rect 2857 2308 2919 2316
rect 2847 2267 2874 2274
rect 2894 2256 2900 2261
rect 2866 2248 2900 2256
rect 2854 2240 2861 2248
rect 2697 2224 2705 2239
rect 2787 2234 2861 2240
rect 2787 2232 2793 2234
rect 2854 2228 2861 2234
rect 2747 2210 2758 2218
rect 2751 2204 2758 2210
rect 2808 2216 2829 2223
rect 2913 2224 2919 2308
rect 2979 2281 2987 2316
rect 3079 2281 3087 2316
rect 3173 2281 3181 2316
rect 2973 2245 2981 2267
rect 3073 2245 3081 2267
rect 3179 2245 3187 2267
rect 3237 2253 3245 2316
rect 3259 2304 3273 2312
rect 3293 2312 3333 2318
rect 3253 2253 3267 2267
rect 2955 2238 2980 2245
rect 3055 2238 3080 2245
rect 3180 2238 3205 2245
rect 2955 2224 2963 2238
rect 2808 2204 2815 2216
rect 2873 2204 2880 2210
rect 2867 2198 2880 2204
rect 2971 2224 3023 2227
rect 3055 2224 3063 2238
rect 2983 2218 3011 2224
rect 3071 2224 3123 2227
rect 3083 2218 3111 2224
rect 3137 2224 3189 2227
rect 3149 2218 3177 2224
rect 3197 2224 3205 2238
rect 3237 2239 3253 2253
rect 3327 2240 3333 2312
rect 3341 2312 3347 2326
rect 3365 2322 3403 2330
rect 3719 2317 3723 2326
rect 3341 2306 3385 2312
rect 3397 2308 3459 2316
rect 3387 2267 3414 2274
rect 3434 2256 3440 2261
rect 3406 2248 3440 2256
rect 3394 2240 3401 2248
rect 3237 2224 3245 2239
rect 3327 2234 3401 2240
rect 3327 2232 3333 2234
rect 3394 2228 3401 2234
rect 3287 2210 3298 2218
rect 3291 2204 3298 2210
rect 3348 2216 3369 2223
rect 3453 2224 3459 2308
rect 3519 2281 3527 2316
rect 3603 2309 3620 2316
rect 3513 2245 3521 2267
rect 3613 2261 3620 2309
rect 3657 2308 3665 2316
rect 3657 2300 3693 2308
rect 3495 2238 3520 2245
rect 3495 2224 3503 2238
rect 3348 2204 3355 2216
rect 3413 2204 3420 2210
rect 3407 2198 3420 2204
rect 3511 2224 3563 2227
rect 3523 2218 3551 2224
rect 3613 2204 3620 2247
rect 3698 2244 3704 2299
rect 3714 2273 3723 2317
rect 3737 2317 3773 2323
rect 3737 2287 3743 2317
rect 3795 2301 3803 2356
rect 3863 2390 3891 2396
rect 3903 2318 3931 2324
rect 3983 2390 4011 2396
rect 4023 2318 4051 2324
rect 4137 2350 4145 2356
rect 4187 2350 4199 2356
rect 4127 2336 4145 2350
rect 4173 2338 4195 2350
rect 4241 2342 4253 2376
rect 4137 2330 4145 2336
rect 4137 2322 4175 2330
rect 4193 2326 4223 2332
rect 3872 2310 3884 2316
rect 3992 2310 4004 2316
rect 3872 2304 3899 2310
rect 3683 2232 3693 2238
rect 3683 2204 3689 2232
rect 3720 2224 3727 2259
rect 3795 2238 3803 2287
rect 3893 2281 3899 2304
rect 3992 2304 4019 2310
rect 3779 2232 3803 2238
rect 3779 2224 3791 2232
rect 3900 2224 3907 2267
rect 3957 2243 3963 2293
rect 4013 2281 4019 2304
rect 4081 2308 4143 2316
rect 3947 2237 3963 2243
rect 4020 2224 4027 2267
rect 4081 2224 4087 2308
rect 4193 2312 4199 2326
rect 4241 2318 4247 2336
rect 4155 2306 4199 2312
rect 4207 2312 4247 2318
rect 4126 2267 4153 2274
rect 4100 2256 4106 2261
rect 4100 2248 4134 2256
rect 4139 2240 4146 2248
rect 4207 2240 4213 2312
rect 4267 2304 4281 2312
rect 4273 2253 4287 2267
rect 4295 2253 4303 2316
rect 4139 2234 4213 2240
rect 4287 2239 4303 2253
rect 4139 2228 4146 2234
rect 4207 2232 4213 2234
rect 2498 2178 2510 2184
rect 2627 2178 2639 2184
rect 2719 2178 2731 2184
rect 2777 2178 2789 2184
rect 2825 2178 2837 2184
rect 2887 2178 2899 2184
rect 2991 2178 3003 2184
rect 3091 2178 3103 2184
rect 3157 2178 3169 2184
rect 3259 2178 3271 2184
rect 3317 2178 3329 2184
rect 3365 2178 3377 2184
rect 3427 2178 3439 2184
rect 3531 2178 3543 2184
rect 3591 2178 3603 2184
rect 3631 2178 3643 2184
rect 3657 2178 3665 2184
rect 3697 2178 3709 2184
rect 3809 2178 3821 2184
rect 3872 2178 3884 2184
rect 3928 2178 3940 2184
rect 4171 2216 4192 2223
rect 4295 2224 4303 2239
rect 4120 2204 4127 2210
rect 4185 2204 4192 2216
rect 4242 2210 4253 2218
rect 4242 2204 4249 2210
rect 4120 2198 4133 2204
rect 4367 2342 4379 2376
rect 4421 2350 4433 2356
rect 4475 2350 4483 2356
rect 4425 2338 4447 2350
rect 4475 2336 4493 2350
rect 4373 2318 4379 2336
rect 4397 2326 4427 2332
rect 4475 2330 4483 2336
rect 4317 2253 4325 2316
rect 4339 2304 4353 2312
rect 4373 2312 4413 2318
rect 4333 2253 4347 2267
rect 4317 2239 4333 2253
rect 4407 2240 4413 2312
rect 4421 2312 4427 2326
rect 4445 2322 4483 2330
rect 4657 2396 4669 2402
rect 4697 2396 4709 2402
rect 4421 2306 4465 2312
rect 4477 2308 4539 2316
rect 4467 2267 4494 2274
rect 4514 2256 4520 2261
rect 4486 2248 4520 2256
rect 4474 2240 4481 2248
rect 4317 2224 4325 2239
rect 4407 2234 4481 2240
rect 4407 2232 4413 2234
rect 4474 2228 4481 2234
rect 4367 2210 4378 2218
rect 4371 2204 4378 2210
rect 4428 2216 4449 2223
rect 4533 2224 4539 2308
rect 4593 2281 4601 2316
rect 4677 2301 4685 2356
rect 4599 2245 4607 2267
rect 4600 2238 4625 2245
rect 4428 2204 4435 2216
rect 4493 2204 4500 2210
rect 4487 2198 4500 2204
rect 4557 2224 4609 2227
rect 4569 2218 4597 2224
rect 4617 2224 4625 2238
rect 4677 2238 4685 2287
rect 4677 2232 4701 2238
rect 4689 2224 4701 2232
rect 3992 2178 4004 2184
rect 4048 2178 4060 2184
rect 4101 2178 4113 2184
rect 4163 2178 4175 2184
rect 4211 2178 4223 2184
rect 4269 2178 4281 2184
rect 4339 2178 4351 2184
rect 4397 2178 4409 2184
rect 4445 2178 4457 2184
rect 4507 2178 4519 2184
rect 4577 2178 4589 2184
rect 4659 2178 4671 2184
rect 4782 2178 4842 2642
rect 4 2176 4842 2178
rect 4776 2164 4842 2176
rect 4 2162 4842 2164
rect 49 2156 61 2162
rect 151 2156 163 2162
rect 270 2156 282 2162
rect 31 2073 39 2116
rect 71 2110 79 2136
rect 57 2104 79 2110
rect 57 2098 60 2104
rect 31 2059 33 2073
rect 31 2024 39 2059
rect 53 2042 60 2098
rect 115 2102 123 2116
rect 143 2116 171 2122
rect 131 2113 183 2116
rect 115 2095 140 2102
rect 216 2098 234 2100
rect 97 2077 113 2083
rect 57 2036 60 2042
rect 57 2030 83 2036
rect 75 1984 83 2030
rect 97 2003 103 2077
rect 133 2073 141 2095
rect 216 2089 246 2098
rect 300 2156 312 2162
rect 350 2156 362 2162
rect 400 2156 412 2162
rect 450 2156 462 2162
rect 340 2116 366 2127
rect 498 2156 510 2162
rect 598 2156 610 2162
rect 700 2156 712 2162
rect 750 2156 762 2162
rect 851 2156 863 2162
rect 898 2156 910 2162
rect 998 2156 1010 2162
rect 1098 2156 1110 2162
rect 1200 2156 1212 2162
rect 1250 2156 1262 2162
rect 440 2116 466 2127
rect 216 2061 224 2089
rect 358 2073 366 2116
rect 139 2024 147 2059
rect 458 2073 466 2116
rect 546 2098 564 2100
rect 534 2089 564 2098
rect 740 2116 766 2127
rect 646 2098 664 2100
rect 634 2089 664 2098
rect 556 2061 564 2089
rect 656 2061 664 2089
rect 758 2073 766 2116
rect 815 2102 823 2116
rect 843 2116 871 2122
rect 831 2113 883 2116
rect 815 2095 840 2102
rect 946 2098 964 2100
rect 833 2073 841 2095
rect 934 2089 964 2098
rect 1046 2098 1064 2100
rect 1034 2089 1064 2098
rect 1297 2156 1309 2162
rect 1337 2156 1349 2162
rect 1429 2156 1441 2162
rect 1509 2156 1521 2162
rect 1240 2116 1266 2127
rect 1146 2098 1164 2100
rect 1134 2089 1164 2098
rect 97 1997 113 2003
rect 215 1992 222 2047
rect 358 2024 366 2059
rect 458 2024 466 2059
rect 297 2018 337 2024
rect 297 2016 309 2018
rect 215 1986 262 1992
rect 215 1984 223 1986
rect 251 1984 262 1986
rect 397 2018 437 2024
rect 397 2016 409 2018
rect 558 1992 565 2047
rect 956 2061 964 2089
rect 1056 2061 1064 2089
rect 1087 2077 1113 2083
rect 1156 2061 1164 2089
rect 1258 2073 1266 2116
rect 1277 2097 1293 2103
rect 658 1992 665 2047
rect 758 2024 766 2059
rect 839 2024 847 2059
rect 518 1986 565 1992
rect 518 1984 529 1986
rect 557 1984 565 1986
rect 618 1986 665 1992
rect 618 1984 629 1986
rect 657 1984 665 1986
rect 697 2018 737 2024
rect 697 2016 709 2018
rect 958 1992 965 2047
rect 1058 1992 1065 2047
rect 1158 1992 1165 2047
rect 1258 2024 1266 2059
rect 1277 2047 1283 2097
rect 1320 2093 1327 2136
rect 1539 2156 1551 2162
rect 1671 2156 1683 2162
rect 1720 2156 1732 2162
rect 1770 2156 1782 2162
rect 1399 2108 1411 2116
rect 1479 2108 1491 2116
rect 1569 2108 1581 2116
rect 1399 2102 1423 2108
rect 1320 2031 1327 2079
rect 1320 2024 1337 2031
rect 918 1986 965 1992
rect 918 1984 929 1986
rect 49 1938 61 1944
rect 116 1938 128 1944
rect 166 1938 178 1944
rect 231 1938 243 1944
rect 271 1938 283 1944
rect 317 1938 329 1944
rect 417 1938 429 1944
rect 497 1938 509 1944
rect 537 1938 549 1944
rect 597 1938 609 1944
rect 637 1938 649 1944
rect 717 1938 729 1944
rect 816 1938 828 1944
rect 866 1938 878 1944
rect 957 1984 965 1986
rect 1018 1986 1065 1992
rect 1018 1984 1029 1986
rect 1057 1984 1065 1986
rect 1118 1986 1165 1992
rect 1118 1984 1129 1986
rect 1157 1984 1165 1986
rect 1197 2018 1237 2024
rect 1197 2016 1209 2018
rect 1377 2023 1383 2053
rect 1415 2053 1423 2102
rect 1447 2097 1463 2103
rect 1479 2102 1503 2108
rect 1367 2017 1383 2023
rect 1415 1984 1423 2039
rect 1457 2023 1463 2097
rect 1495 2053 1503 2102
rect 1557 2102 1581 2108
rect 1635 2102 1643 2116
rect 1663 2116 1691 2122
rect 1817 2156 1829 2162
rect 1857 2156 1869 2162
rect 1951 2156 1963 2162
rect 2017 2156 2029 2162
rect 2151 2156 2163 2162
rect 2211 2156 2223 2162
rect 2251 2156 2263 2162
rect 2291 2156 2303 2162
rect 2331 2156 2343 2162
rect 2371 2156 2383 2162
rect 1760 2116 1786 2127
rect 1651 2113 1703 2116
rect 1557 2053 1565 2102
rect 1635 2095 1660 2102
rect 1653 2073 1661 2095
rect 1778 2073 1786 2116
rect 1840 2093 1847 2136
rect 1915 2102 1923 2116
rect 1943 2116 1971 2122
rect 1931 2113 1983 2116
rect 2009 2116 2037 2122
rect 1997 2113 2049 2116
rect 2057 2102 2065 2116
rect 1915 2095 1940 2102
rect 2040 2095 2065 2102
rect 2115 2102 2123 2116
rect 2143 2116 2171 2122
rect 2399 2156 2411 2162
rect 2521 2156 2533 2162
rect 2577 2156 2585 2162
rect 2617 2156 2629 2162
rect 2729 2156 2741 2162
rect 2131 2113 2183 2116
rect 2232 2110 2244 2116
rect 2272 2110 2284 2116
rect 2311 2110 2323 2116
rect 2352 2110 2364 2116
rect 2226 2109 2244 2110
rect 2225 2102 2244 2109
rect 2258 2102 2284 2110
rect 2298 2102 2323 2110
rect 2337 2102 2364 2110
rect 2429 2108 2441 2116
rect 2417 2102 2441 2108
rect 2491 2116 2501 2126
rect 2115 2095 2140 2102
rect 1457 2017 1473 2023
rect 1495 1984 1503 2039
rect 1557 1984 1565 2039
rect 1659 2024 1667 2059
rect 1778 2024 1786 2059
rect 1840 2031 1847 2079
rect 1933 2073 1941 2095
rect 2039 2073 2047 2095
rect 2133 2073 2141 2095
rect 2225 2081 2232 2102
rect 2258 2096 2266 2102
rect 2298 2096 2306 2102
rect 2337 2096 2345 2102
rect 2250 2084 2266 2096
rect 2290 2084 2306 2096
rect 2330 2084 2345 2096
rect 2227 2067 2232 2081
rect 1840 2024 1857 2031
rect 1939 2024 1947 2059
rect 2033 2024 2041 2059
rect 2139 2024 2147 2059
rect 2225 2038 2232 2067
rect 2258 2038 2266 2084
rect 2298 2038 2306 2084
rect 2337 2038 2345 2084
rect 2417 2053 2425 2102
rect 2491 2073 2499 2116
rect 2551 2106 2563 2116
rect 2525 2098 2563 2106
rect 2603 2108 2609 2136
rect 2759 2156 2771 2162
rect 2861 2156 2873 2162
rect 2923 2156 2935 2162
rect 2971 2156 2983 2162
rect 3029 2156 3041 2162
rect 3098 2156 3110 2162
rect 3148 2156 3160 2162
rect 2603 2102 2613 2108
rect 2491 2059 2493 2073
rect 2225 2030 2243 2038
rect 2258 2030 2283 2038
rect 2298 2030 2323 2038
rect 2337 2030 2363 2038
rect 2231 2024 2243 2030
rect 2271 2024 2283 2030
rect 2311 2024 2323 2030
rect 2351 2024 2363 2030
rect 897 1938 909 1944
rect 937 1938 949 1944
rect 997 1938 1009 1944
rect 1037 1938 1049 1944
rect 1097 1938 1109 1944
rect 1137 1938 1149 1944
rect 1217 1938 1229 1944
rect 1297 1938 1309 1944
rect 1391 1938 1403 1944
rect 1431 1938 1443 1944
rect 1471 1938 1483 1944
rect 1511 1938 1523 1944
rect 1537 1938 1549 1944
rect 1577 1938 1589 1944
rect 1717 2018 1757 2024
rect 1717 2016 1729 2018
rect 1636 1938 1648 1944
rect 1686 1938 1698 1944
rect 1737 1938 1749 1944
rect 1817 1938 1829 1944
rect 1916 1938 1928 1944
rect 1966 1938 1978 1944
rect 2002 1938 2014 1944
rect 2052 1938 2064 1944
rect 2116 1938 2128 1944
rect 2166 1938 2178 1944
rect 2417 1984 2425 2039
rect 2491 2024 2499 2059
rect 2211 1938 2223 1944
rect 2251 1938 2263 1944
rect 2291 1938 2303 1944
rect 2331 1938 2343 1944
rect 2371 1938 2383 1944
rect 2534 1984 2542 2098
rect 2618 2041 2624 2096
rect 2640 2081 2647 2116
rect 2699 2108 2711 2116
rect 2789 2108 2801 2116
rect 2699 2102 2723 2108
rect 2577 2032 2613 2040
rect 2577 2024 2585 2032
rect 2634 2023 2643 2067
rect 2715 2053 2723 2102
rect 2777 2102 2801 2108
rect 2880 2136 2893 2142
rect 2880 2130 2887 2136
rect 2945 2124 2952 2136
rect 2777 2053 2785 2102
rect 2639 2014 2643 2023
rect 2715 1984 2723 2039
rect 2777 1984 2785 2039
rect 2841 2032 2847 2116
rect 2931 2117 2952 2124
rect 3002 2130 3009 2136
rect 3002 2122 3013 2130
rect 2899 2106 2906 2112
rect 2967 2106 2973 2108
rect 2899 2100 2973 2106
rect 3055 2101 3063 2116
rect 2899 2092 2906 2100
rect 2860 2084 2894 2092
rect 2860 2079 2866 2084
rect 2886 2066 2913 2073
rect 2841 2024 2903 2032
rect 2915 2028 2959 2034
rect 2397 1938 2409 1944
rect 2437 1938 2449 1944
rect 2507 1938 2519 1944
rect 2551 1938 2563 1944
rect 2607 1938 2619 1944
rect 2691 1938 2703 1944
rect 2731 1938 2743 1944
rect 2897 2010 2935 2018
rect 2953 2014 2959 2028
rect 2967 2028 2973 2100
rect 3047 2087 3063 2101
rect 3033 2073 3047 2087
rect 2967 2022 3007 2028
rect 3027 2028 3041 2036
rect 3055 2024 3063 2087
rect 3094 2116 3120 2127
rect 3177 2156 3189 2162
rect 3217 2156 3229 2162
rect 3292 2156 3304 2162
rect 3348 2156 3360 2162
rect 3401 2156 3413 2162
rect 3463 2156 3475 2162
rect 3511 2156 3523 2162
rect 3569 2156 3581 2162
rect 3637 2156 3649 2162
rect 3741 2156 3753 2162
rect 3803 2156 3815 2162
rect 3851 2156 3863 2162
rect 3909 2156 3921 2162
rect 3979 2156 3991 2162
rect 4037 2156 4049 2162
rect 4085 2156 4097 2162
rect 4147 2156 4159 2162
rect 4232 2156 4244 2162
rect 4288 2156 4300 2162
rect 3094 2073 3102 2116
rect 3200 2093 3207 2136
rect 3420 2136 3433 2142
rect 3420 2130 3427 2136
rect 3485 2124 3492 2136
rect 3094 2024 3102 2059
rect 3200 2031 3207 2079
rect 3320 2073 3327 2116
rect 3313 2036 3319 2059
rect 3200 2024 3217 2031
rect 3292 2030 3319 2036
rect 3381 2032 3387 2116
rect 3471 2117 3492 2124
rect 3542 2130 3549 2136
rect 3542 2122 3553 2130
rect 3439 2106 3446 2112
rect 3507 2106 3513 2108
rect 3439 2100 3513 2106
rect 3595 2101 3603 2116
rect 3629 2116 3657 2122
rect 3617 2113 3669 2116
rect 3760 2136 3773 2142
rect 3760 2130 3767 2136
rect 3825 2124 3832 2136
rect 3677 2102 3685 2116
rect 3439 2092 3446 2100
rect 3400 2084 3434 2092
rect 3400 2079 3406 2084
rect 3426 2066 3453 2073
rect 3292 2024 3304 2030
rect 3381 2024 3443 2032
rect 3455 2028 3499 2034
rect 2897 2004 2905 2010
rect 2953 2008 2983 2014
rect 3001 2004 3007 2022
rect 2887 1990 2905 2004
rect 2933 1990 2955 2002
rect 2897 1984 2905 1990
rect 2947 1984 2959 1990
rect 3001 1964 3013 1998
rect 3123 2018 3163 2024
rect 3151 2016 3163 2018
rect 3283 1944 3311 1950
rect 3323 2016 3351 2022
rect 3437 2010 3475 2018
rect 3493 2014 3499 2028
rect 3507 2028 3513 2100
rect 3587 2087 3603 2101
rect 3660 2095 3685 2102
rect 3573 2073 3587 2087
rect 3507 2022 3547 2028
rect 3567 2028 3581 2036
rect 3595 2024 3603 2087
rect 3659 2073 3667 2095
rect 3653 2024 3661 2059
rect 3721 2032 3727 2116
rect 3811 2117 3832 2124
rect 3882 2130 3889 2136
rect 3882 2122 3893 2130
rect 3779 2106 3786 2112
rect 3847 2106 3853 2108
rect 3779 2100 3853 2106
rect 3935 2101 3943 2116
rect 3779 2092 3786 2100
rect 3740 2084 3774 2092
rect 3740 2079 3746 2084
rect 3766 2066 3793 2073
rect 3721 2024 3783 2032
rect 3795 2028 3839 2034
rect 3437 2004 3445 2010
rect 3493 2008 3523 2014
rect 3541 2004 3547 2022
rect 3427 1990 3445 2004
rect 3473 1990 3495 2002
rect 3437 1984 3445 1990
rect 3487 1984 3499 1990
rect 3541 1964 3553 1998
rect 3777 2010 3815 2018
rect 3833 2014 3839 2028
rect 3847 2028 3853 2100
rect 3927 2087 3943 2101
rect 3913 2073 3927 2087
rect 3847 2022 3887 2028
rect 3907 2028 3921 2036
rect 3935 2024 3943 2087
rect 3777 2004 3785 2010
rect 3833 2008 3863 2014
rect 3881 2004 3887 2022
rect 3767 1990 3785 2004
rect 3813 1990 3835 2002
rect 3777 1984 3785 1990
rect 3827 1984 3839 1990
rect 3881 1964 3893 1998
rect 4127 2136 4140 2142
rect 4011 2130 4018 2136
rect 4007 2122 4018 2130
rect 4068 2124 4075 2136
rect 4133 2130 4140 2136
rect 3957 2101 3965 2116
rect 4068 2117 4089 2124
rect 4317 2156 4329 2162
rect 4391 2156 4403 2162
rect 4431 2156 4443 2162
rect 4471 2156 4483 2162
rect 4511 2156 4523 2162
rect 4559 2156 4571 2162
rect 4617 2156 4629 2162
rect 4665 2156 4677 2162
rect 4727 2156 4739 2162
rect 4047 2106 4053 2108
rect 4114 2106 4121 2112
rect 3957 2087 3973 2101
rect 4047 2100 4121 2106
rect 3957 2024 3965 2087
rect 3973 2073 3987 2087
rect 3979 2028 3993 2036
rect 4047 2028 4053 2100
rect 4114 2092 4121 2100
rect 4126 2084 4160 2092
rect 4154 2079 4160 2084
rect 4107 2066 4134 2073
rect 4013 2022 4053 2028
rect 4061 2028 4105 2034
rect 4013 2004 4019 2022
rect 4061 2014 4067 2028
rect 4173 2032 4179 2116
rect 4260 2073 4267 2116
rect 4336 2081 4344 2136
rect 4413 2093 4420 2136
rect 4493 2093 4500 2136
rect 4707 2136 4720 2142
rect 4591 2130 4598 2136
rect 4587 2122 4598 2130
rect 4648 2124 4655 2136
rect 4713 2130 4720 2136
rect 4537 2101 4545 2116
rect 4648 2117 4669 2124
rect 4627 2106 4633 2108
rect 4694 2106 4701 2112
rect 4537 2087 4553 2101
rect 4627 2100 4701 2106
rect 4253 2036 4259 2059
rect 4117 2024 4179 2032
rect 4232 2030 4259 2036
rect 4232 2024 4244 2030
rect 4037 2008 4067 2014
rect 4085 2010 4123 2018
rect 4115 2004 4123 2010
rect 4007 1964 4019 1998
rect 4065 1990 4087 2002
rect 4115 1990 4133 2004
rect 4061 1984 4073 1990
rect 4115 1984 4123 1990
rect 4223 1944 4251 1950
rect 4263 2016 4291 2022
rect 4336 1984 4344 2067
rect 4413 2031 4420 2079
rect 4493 2031 4500 2079
rect 4403 2024 4420 2031
rect 4483 2024 4500 2031
rect 4537 2024 4545 2087
rect 4553 2073 4567 2087
rect 4559 2028 4573 2036
rect 4627 2028 4633 2100
rect 4694 2092 4701 2100
rect 4706 2084 4740 2092
rect 4734 2079 4740 2084
rect 4687 2066 4714 2073
rect 4593 2022 4633 2028
rect 4641 2028 4685 2034
rect 4593 2004 4599 2022
rect 4641 2014 4647 2028
rect 4753 2032 4759 2116
rect 4697 2024 4759 2032
rect 4617 2008 4647 2014
rect 4665 2010 4703 2018
rect 4695 2004 4703 2010
rect 4587 1964 4599 1998
rect 4645 1990 4667 2002
rect 4695 1990 4713 2004
rect 4641 1984 4653 1990
rect 4695 1984 4703 1990
rect 2757 1938 2769 1944
rect 2797 1938 2809 1944
rect 2861 1938 2873 1944
rect 2927 1938 2939 1944
rect 2973 1938 2985 1944
rect 3031 1938 3043 1944
rect 3131 1938 3143 1944
rect 3177 1938 3189 1944
rect 3331 1938 3343 1944
rect 3401 1938 3413 1944
rect 3467 1938 3479 1944
rect 3513 1938 3525 1944
rect 3571 1938 3583 1944
rect 3622 1938 3634 1944
rect 3672 1938 3684 1944
rect 3741 1938 3753 1944
rect 3807 1938 3819 1944
rect 3853 1938 3865 1944
rect 3911 1938 3923 1944
rect 3977 1938 3989 1944
rect 4035 1938 4047 1944
rect 4081 1938 4093 1944
rect 4147 1938 4159 1944
rect 4271 1938 4283 1944
rect 4317 1938 4329 1944
rect 4431 1938 4443 1944
rect 4511 1938 4523 1944
rect 4557 1938 4569 1944
rect 4615 1938 4627 1944
rect 4661 1938 4673 1944
rect 4727 1938 4739 1944
rect -62 1936 4776 1938
rect -62 1924 4 1936
rect -62 1922 4776 1924
rect -62 1458 -2 1922
rect 91 1916 103 1922
rect 142 1916 154 1922
rect 192 1916 204 1922
rect 43 1910 71 1916
rect 83 1838 111 1844
rect 237 1916 249 1922
rect 277 1916 289 1922
rect 351 1916 363 1922
rect 391 1916 403 1922
rect 437 1916 449 1922
rect 537 1916 549 1922
rect 581 1916 593 1922
rect 671 1916 683 1922
rect 719 1916 731 1922
rect 796 1916 808 1922
rect 846 1916 858 1922
rect 52 1830 64 1836
rect 52 1824 79 1830
rect 73 1801 79 1824
rect 173 1801 181 1836
rect 80 1744 87 1787
rect 179 1765 187 1787
rect 217 1783 223 1833
rect 257 1821 265 1876
rect 335 1874 343 1876
rect 371 1874 382 1876
rect 335 1868 382 1874
rect 335 1813 342 1868
rect 429 1838 457 1844
rect 469 1910 497 1916
rect 476 1830 488 1836
rect 461 1824 488 1830
rect 207 1777 223 1783
rect 180 1758 205 1765
rect 137 1744 189 1747
rect 149 1738 177 1744
rect 197 1744 205 1758
rect 257 1758 265 1807
rect 461 1801 467 1824
rect 336 1771 344 1799
rect 336 1762 366 1771
rect 336 1760 354 1762
rect 257 1752 281 1758
rect 269 1744 281 1752
rect 453 1744 460 1787
rect 558 1762 566 1876
rect 601 1801 609 1836
rect 656 1801 664 1836
rect 697 1830 705 1876
rect 882 1916 894 1922
rect 932 1916 944 1922
rect 977 1916 989 1922
rect 1017 1916 1029 1922
rect 1077 1916 1089 1922
rect 1137 1916 1149 1922
rect 1177 1916 1189 1922
rect 1237 1916 1249 1922
rect 1277 1916 1289 1922
rect 1371 1916 1383 1922
rect 1471 1916 1483 1922
rect 1517 1916 1529 1922
rect 1557 1916 1569 1922
rect 1617 1916 1629 1922
rect 1711 1916 1723 1922
rect 1771 1916 1783 1922
rect 1811 1916 1823 1922
rect 998 1874 1009 1876
rect 1037 1874 1045 1876
rect 998 1868 1045 1874
rect 697 1824 723 1830
rect 720 1818 723 1824
rect 607 1787 609 1801
rect 537 1754 575 1762
rect 537 1744 549 1754
rect 601 1744 609 1787
rect 656 1744 664 1787
rect 720 1762 727 1818
rect 741 1801 749 1836
rect 819 1801 827 1836
rect 913 1801 921 1836
rect 1038 1813 1045 1868
rect 747 1787 749 1801
rect 720 1756 723 1762
rect 701 1750 723 1756
rect 52 1698 64 1704
rect 108 1698 120 1704
rect 157 1698 169 1704
rect 239 1698 251 1704
rect 390 1698 402 1704
rect 599 1734 609 1744
rect 701 1724 709 1750
rect 741 1744 749 1787
rect 813 1765 821 1787
rect 919 1765 927 1787
rect 1036 1771 1044 1799
rect 1096 1793 1104 1876
rect 1158 1874 1169 1876
rect 1197 1874 1205 1876
rect 1158 1868 1205 1874
rect 1258 1874 1269 1876
rect 1297 1874 1305 1876
rect 1258 1868 1305 1874
rect 1117 1857 1133 1863
rect 795 1758 820 1765
rect 920 1758 945 1765
rect 795 1744 803 1758
rect 811 1744 863 1747
rect 823 1738 851 1744
rect 877 1744 929 1747
rect 889 1738 917 1744
rect 937 1744 945 1758
rect 1014 1762 1044 1771
rect 1117 1783 1123 1857
rect 1198 1813 1205 1868
rect 1298 1813 1305 1868
rect 1026 1760 1044 1762
rect 1096 1724 1104 1779
rect 1117 1777 1153 1783
rect 1196 1771 1204 1799
rect 1296 1771 1304 1799
rect 1356 1793 1364 1876
rect 1423 1910 1451 1916
rect 1463 1838 1491 1844
rect 1538 1874 1549 1876
rect 1577 1874 1585 1876
rect 1538 1868 1585 1874
rect 1432 1830 1444 1836
rect 1432 1824 1459 1830
rect 1453 1801 1459 1824
rect 1578 1813 1585 1868
rect 1174 1762 1204 1771
rect 1186 1760 1204 1762
rect 1274 1762 1304 1771
rect 1286 1760 1304 1762
rect 1356 1724 1364 1779
rect 1460 1744 1467 1787
rect 1576 1771 1584 1799
rect 1636 1793 1644 1876
rect 1755 1874 1763 1876
rect 1837 1916 1849 1922
rect 1881 1916 1893 1922
rect 1961 1916 1973 1922
rect 2027 1916 2039 1922
rect 2073 1916 2085 1922
rect 2131 1916 2143 1922
rect 2231 1916 2243 1922
rect 1791 1874 1802 1876
rect 1755 1868 1802 1874
rect 1696 1801 1704 1836
rect 1755 1813 1762 1868
rect 420 1698 432 1704
rect 476 1698 488 1704
rect 567 1698 579 1704
rect 671 1698 683 1704
rect 719 1698 731 1704
rect 831 1698 843 1704
rect 897 1698 909 1704
rect 978 1698 990 1704
rect 1077 1698 1089 1704
rect 1138 1698 1150 1704
rect 1238 1698 1250 1704
rect 1371 1698 1383 1704
rect 1432 1698 1444 1704
rect 1488 1698 1500 1704
rect 1554 1762 1584 1771
rect 1566 1760 1584 1762
rect 1636 1724 1644 1779
rect 1696 1744 1704 1787
rect 1756 1771 1764 1799
rect 1756 1762 1786 1771
rect 1756 1760 1774 1762
rect 1858 1762 1866 1876
rect 1997 1870 2005 1876
rect 2047 1870 2059 1876
rect 1987 1856 2005 1870
rect 2033 1858 2055 1870
rect 2101 1862 2113 1896
rect 1997 1850 2005 1856
rect 1997 1842 2035 1850
rect 2053 1846 2083 1852
rect 1901 1801 1909 1836
rect 1907 1787 1909 1801
rect 1837 1754 1875 1762
rect 1837 1744 1849 1754
rect 1901 1744 1909 1787
rect 1899 1734 1909 1744
rect 1941 1828 2003 1836
rect 1941 1744 1947 1828
rect 2053 1832 2059 1846
rect 2101 1838 2107 1856
rect 2015 1826 2059 1832
rect 2067 1832 2107 1838
rect 1986 1787 2013 1794
rect 1960 1776 1966 1781
rect 1960 1768 1994 1776
rect 1999 1760 2006 1768
rect 2067 1760 2073 1832
rect 2127 1824 2141 1832
rect 2133 1773 2147 1787
rect 2155 1773 2163 1836
rect 2257 1916 2269 1922
rect 2322 1916 2334 1922
rect 2372 1916 2384 1922
rect 2203 1829 2220 1836
rect 1999 1754 2073 1760
rect 2147 1759 2163 1773
rect 1999 1748 2006 1754
rect 2067 1752 2073 1754
rect 2031 1736 2052 1743
rect 2155 1744 2163 1759
rect 1980 1724 1987 1730
rect 2045 1724 2052 1736
rect 2102 1730 2113 1738
rect 2102 1724 2109 1730
rect 1980 1718 1993 1724
rect 2213 1781 2220 1829
rect 2276 1793 2284 1876
rect 2417 1916 2429 1922
rect 2497 1916 2509 1922
rect 2582 1916 2594 1922
rect 2632 1916 2644 1922
rect 2691 1916 2703 1922
rect 2731 1916 2743 1922
rect 2811 1916 2823 1922
rect 2353 1801 2361 1836
rect 2440 1829 2457 1836
rect 2520 1829 2537 1836
rect 2213 1724 2220 1767
rect 2276 1724 2284 1779
rect 2359 1765 2367 1787
rect 2440 1781 2447 1829
rect 2520 1781 2527 1829
rect 2613 1801 2621 1836
rect 2715 1821 2723 1876
rect 2842 1916 2854 1922
rect 2892 1916 2904 1922
rect 2937 1916 2949 1922
rect 3051 1916 3063 1922
rect 3097 1916 3109 1922
rect 3155 1916 3167 1922
rect 3201 1916 3213 1922
rect 3267 1916 3279 1922
rect 3322 1916 3334 1922
rect 3372 1916 3384 1922
rect 2783 1829 2800 1836
rect 2360 1758 2385 1765
rect 2317 1744 2369 1747
rect 1518 1698 1530 1704
rect 1617 1698 1629 1704
rect 1711 1698 1723 1704
rect 1810 1698 1822 1704
rect 1867 1698 1879 1704
rect 1961 1698 1973 1704
rect 2023 1698 2035 1704
rect 2071 1698 2083 1704
rect 2129 1698 2141 1704
rect 2191 1698 2203 1704
rect 2231 1698 2243 1704
rect 2329 1738 2357 1744
rect 2377 1744 2385 1758
rect 2440 1724 2447 1767
rect 2520 1724 2527 1767
rect 2619 1765 2627 1787
rect 2620 1758 2645 1765
rect 2715 1758 2723 1807
rect 2577 1744 2629 1747
rect 2257 1698 2269 1704
rect 2337 1698 2349 1704
rect 2417 1698 2429 1704
rect 2457 1698 2469 1704
rect 2589 1738 2617 1744
rect 2637 1744 2645 1758
rect 2699 1752 2723 1758
rect 2793 1781 2800 1829
rect 2873 1801 2881 1836
rect 2956 1793 2964 1876
rect 3127 1862 3139 1896
rect 3181 1870 3193 1876
rect 3235 1870 3243 1876
rect 3185 1858 3207 1870
rect 3235 1856 3253 1870
rect 3133 1838 3139 1856
rect 3157 1846 3187 1852
rect 3235 1850 3243 1856
rect 3023 1829 3040 1836
rect 2699 1744 2711 1752
rect 2793 1724 2800 1767
rect 2879 1765 2887 1787
rect 3033 1781 3040 1829
rect 2880 1758 2905 1765
rect 2837 1744 2889 1747
rect 2497 1698 2509 1704
rect 2537 1698 2549 1704
rect 2597 1698 2609 1704
rect 2729 1698 2741 1704
rect 2849 1738 2877 1744
rect 2897 1744 2905 1758
rect 2956 1724 2964 1779
rect 3077 1773 3085 1836
rect 3099 1824 3113 1832
rect 3133 1832 3173 1838
rect 3093 1773 3107 1787
rect 3033 1724 3040 1767
rect 3077 1759 3093 1773
rect 3167 1760 3173 1832
rect 3181 1832 3187 1846
rect 3205 1842 3243 1850
rect 3417 1916 3429 1922
rect 3457 1916 3469 1922
rect 3517 1916 3529 1922
rect 3575 1916 3587 1922
rect 3621 1916 3633 1922
rect 3687 1916 3699 1922
rect 3759 1916 3771 1922
rect 3831 1916 3843 1922
rect 3871 1916 3883 1922
rect 3181 1826 3225 1832
rect 3237 1828 3299 1836
rect 3227 1787 3254 1794
rect 3274 1776 3280 1781
rect 3246 1768 3280 1776
rect 3234 1760 3241 1768
rect 3077 1744 3085 1759
rect 3167 1754 3241 1760
rect 3167 1752 3173 1754
rect 3234 1748 3241 1754
rect 3127 1730 3138 1738
rect 3131 1724 3138 1730
rect 3188 1736 3209 1743
rect 3293 1744 3299 1828
rect 3353 1801 3361 1836
rect 3437 1821 3445 1876
rect 3547 1862 3559 1896
rect 3601 1870 3613 1876
rect 3655 1870 3663 1876
rect 3605 1858 3627 1870
rect 3655 1856 3673 1870
rect 3553 1838 3559 1856
rect 3577 1846 3607 1852
rect 3655 1850 3663 1856
rect 3359 1765 3367 1787
rect 3360 1758 3385 1765
rect 3188 1724 3195 1736
rect 3253 1724 3260 1730
rect 3247 1718 3260 1724
rect 3317 1744 3369 1747
rect 3329 1738 3357 1744
rect 3377 1744 3385 1758
rect 3437 1758 3445 1807
rect 3497 1773 3505 1836
rect 3519 1824 3533 1832
rect 3553 1832 3593 1838
rect 3513 1773 3527 1787
rect 3497 1759 3513 1773
rect 3587 1760 3593 1832
rect 3601 1832 3607 1846
rect 3625 1842 3663 1850
rect 3601 1826 3645 1832
rect 3657 1828 3719 1836
rect 3647 1787 3674 1794
rect 3694 1776 3700 1781
rect 3666 1768 3700 1776
rect 3654 1760 3661 1768
rect 3437 1752 3461 1758
rect 3449 1744 3461 1752
rect 3497 1744 3505 1759
rect 3587 1754 3661 1760
rect 3587 1752 3593 1754
rect 3654 1748 3661 1754
rect 3547 1730 3558 1738
rect 3551 1724 3558 1730
rect 3608 1736 3629 1743
rect 3713 1744 3719 1828
rect 3737 1830 3745 1876
rect 3916 1916 3928 1922
rect 3966 1916 3978 1922
rect 3737 1824 3763 1830
rect 3760 1818 3763 1824
rect 3760 1762 3767 1818
rect 3781 1801 3789 1836
rect 3855 1821 3863 1876
rect 3897 1857 3913 1863
rect 3787 1787 3789 1801
rect 3760 1756 3763 1762
rect 3608 1724 3615 1736
rect 3673 1724 3680 1730
rect 3667 1718 3680 1724
rect 3741 1750 3763 1756
rect 3741 1724 3749 1750
rect 3781 1744 3789 1787
rect 3855 1758 3863 1807
rect 3897 1783 3903 1857
rect 4016 1916 4028 1922
rect 4066 1916 4078 1922
rect 4127 1916 4139 1922
rect 4231 1916 4243 1922
rect 4277 1916 4289 1922
rect 4411 1916 4423 1922
rect 4457 1916 4469 1922
rect 4515 1916 4527 1922
rect 4561 1916 4573 1922
rect 4627 1916 4639 1922
rect 4691 1916 4703 1922
rect 4731 1916 4743 1922
rect 4159 1837 4163 1846
rect 3939 1801 3947 1836
rect 4039 1801 4047 1836
rect 4097 1828 4105 1836
rect 4097 1820 4133 1828
rect 3897 1777 3913 1783
rect 3933 1765 3941 1787
rect 4033 1765 4041 1787
rect 3839 1752 3863 1758
rect 3915 1758 3940 1765
rect 4015 1758 4040 1765
rect 4138 1764 4144 1819
rect 4154 1793 4163 1837
rect 4216 1793 4224 1876
rect 4257 1842 4269 1844
rect 4257 1836 4297 1842
rect 4487 1862 4499 1896
rect 4541 1870 4553 1876
rect 4595 1870 4603 1876
rect 4545 1858 4567 1870
rect 4595 1856 4613 1870
rect 4493 1838 4499 1856
rect 4517 1846 4547 1852
rect 4595 1850 4603 1856
rect 4318 1801 4326 1836
rect 4383 1829 4400 1836
rect 3839 1744 3851 1752
rect 3915 1744 3923 1758
rect 3931 1744 3983 1747
rect 4015 1744 4023 1758
rect 4123 1752 4133 1758
rect 3943 1738 3971 1744
rect 4031 1744 4083 1747
rect 4043 1738 4071 1744
rect 4123 1724 4129 1752
rect 4160 1744 4167 1779
rect 4216 1724 4224 1779
rect 4318 1744 4326 1787
rect 2771 1698 2783 1704
rect 2811 1698 2823 1704
rect 2857 1698 2869 1704
rect 2937 1698 2949 1704
rect 3011 1698 3023 1704
rect 3051 1698 3063 1704
rect 3099 1698 3111 1704
rect 3157 1698 3169 1704
rect 3205 1698 3217 1704
rect 3267 1698 3279 1704
rect 3337 1698 3349 1704
rect 3419 1698 3431 1704
rect 3519 1698 3531 1704
rect 3577 1698 3589 1704
rect 3625 1698 3637 1704
rect 3687 1698 3699 1704
rect 3759 1698 3771 1704
rect 3869 1698 3881 1704
rect 3951 1698 3963 1704
rect 4051 1698 4063 1704
rect 4097 1698 4105 1704
rect 4137 1698 4149 1704
rect 4231 1698 4243 1704
rect 4300 1733 4326 1744
rect 4393 1781 4400 1829
rect 4437 1773 4445 1836
rect 4459 1824 4473 1832
rect 4493 1832 4533 1838
rect 4453 1773 4467 1787
rect 4393 1724 4400 1767
rect 4437 1759 4453 1773
rect 4527 1760 4533 1832
rect 4541 1832 4547 1846
rect 4565 1842 4603 1850
rect 4541 1826 4585 1832
rect 4597 1828 4659 1836
rect 4587 1787 4614 1794
rect 4634 1776 4640 1781
rect 4606 1768 4640 1776
rect 4594 1760 4601 1768
rect 4437 1744 4445 1759
rect 4527 1754 4601 1760
rect 4527 1752 4533 1754
rect 4260 1698 4272 1704
rect 4310 1698 4322 1704
rect 4594 1748 4601 1754
rect 4487 1730 4498 1738
rect 4491 1724 4498 1730
rect 4548 1736 4569 1743
rect 4653 1744 4659 1828
rect 4715 1821 4723 1876
rect 4715 1758 4723 1807
rect 4548 1724 4555 1736
rect 4613 1724 4620 1730
rect 4607 1718 4620 1724
rect 4699 1752 4723 1758
rect 4699 1744 4711 1752
rect 4371 1698 4383 1704
rect 4411 1698 4423 1704
rect 4459 1698 4471 1704
rect 4517 1698 4529 1704
rect 4565 1698 4577 1704
rect 4627 1698 4639 1704
rect 4729 1698 4741 1704
rect 4782 1698 4842 2162
rect 4 1696 4842 1698
rect 4776 1684 4842 1696
rect 4 1682 4842 1684
rect 51 1676 63 1682
rect 98 1676 110 1682
rect 148 1676 160 1682
rect 36 1601 44 1656
rect 94 1636 120 1647
rect 178 1676 190 1682
rect 279 1676 291 1682
rect 411 1676 423 1682
rect 489 1676 501 1682
rect 571 1676 583 1682
rect 94 1593 102 1636
rect 309 1628 321 1636
rect 226 1618 244 1620
rect 36 1504 44 1587
rect 214 1609 244 1618
rect 236 1581 244 1609
rect 257 1617 273 1623
rect 94 1544 102 1579
rect 123 1538 163 1544
rect 151 1536 163 1538
rect 238 1512 245 1567
rect 257 1543 263 1617
rect 297 1622 321 1628
rect 375 1622 383 1636
rect 403 1636 431 1642
rect 598 1676 610 1682
rect 700 1676 712 1682
rect 750 1676 762 1682
rect 391 1633 443 1636
rect 297 1573 305 1622
rect 375 1615 400 1622
rect 393 1593 401 1615
rect 471 1593 479 1636
rect 511 1630 519 1656
rect 497 1624 519 1630
rect 497 1618 500 1624
rect 471 1579 473 1593
rect 257 1537 273 1543
rect 198 1506 245 1512
rect 198 1504 209 1506
rect 237 1504 245 1506
rect 297 1504 305 1559
rect 399 1544 407 1579
rect 471 1544 479 1579
rect 493 1562 500 1618
rect 556 1601 564 1656
rect 798 1676 810 1682
rect 900 1676 912 1682
rect 950 1676 962 1682
rect 740 1636 766 1647
rect 646 1618 664 1620
rect 634 1609 664 1618
rect 497 1556 500 1562
rect 497 1550 523 1556
rect 51 1458 63 1464
rect 131 1458 143 1464
rect 177 1458 189 1464
rect 217 1458 229 1464
rect 277 1458 289 1464
rect 317 1458 329 1464
rect 515 1504 523 1550
rect 556 1504 564 1587
rect 656 1581 664 1609
rect 758 1593 766 1636
rect 998 1676 1010 1682
rect 1151 1676 1163 1682
rect 1198 1676 1210 1682
rect 1300 1676 1312 1682
rect 1350 1676 1362 1682
rect 1431 1676 1443 1682
rect 940 1636 966 1647
rect 846 1618 864 1620
rect 834 1609 864 1618
rect 856 1581 864 1609
rect 958 1593 966 1636
rect 1046 1618 1064 1620
rect 1034 1609 1064 1618
rect 1115 1622 1123 1636
rect 1143 1636 1171 1642
rect 1131 1633 1183 1636
rect 1115 1615 1140 1622
rect 1267 1637 1283 1643
rect 1246 1618 1264 1620
rect 658 1512 665 1567
rect 758 1544 766 1579
rect 1056 1581 1064 1609
rect 618 1506 665 1512
rect 618 1504 629 1506
rect 376 1458 388 1464
rect 426 1458 438 1464
rect 489 1458 501 1464
rect 571 1458 583 1464
rect 657 1504 665 1506
rect 697 1538 737 1544
rect 697 1536 709 1538
rect 858 1512 865 1567
rect 958 1544 966 1579
rect 818 1506 865 1512
rect 818 1504 829 1506
rect 857 1504 865 1506
rect 897 1538 937 1544
rect 897 1536 909 1538
rect 1058 1512 1065 1567
rect 1077 1543 1083 1613
rect 1133 1593 1141 1615
rect 1234 1609 1264 1618
rect 1256 1581 1264 1609
rect 1077 1537 1093 1543
rect 1139 1544 1147 1579
rect 1018 1506 1065 1512
rect 1018 1504 1029 1506
rect 1057 1504 1065 1506
rect 1258 1512 1265 1567
rect 1277 1563 1283 1637
rect 1458 1676 1470 1682
rect 1560 1676 1572 1682
rect 1610 1676 1622 1682
rect 1340 1636 1366 1647
rect 1358 1593 1366 1636
rect 1416 1601 1424 1656
rect 1658 1676 1670 1682
rect 1777 1676 1789 1682
rect 1878 1676 1890 1682
rect 1928 1676 1940 1682
rect 1600 1636 1626 1647
rect 1506 1618 1524 1620
rect 1494 1609 1524 1618
rect 1277 1557 1293 1563
rect 1358 1544 1366 1579
rect 1218 1506 1265 1512
rect 1218 1504 1229 1506
rect 597 1458 609 1464
rect 637 1458 649 1464
rect 717 1458 729 1464
rect 797 1458 809 1464
rect 837 1458 849 1464
rect 917 1458 929 1464
rect 997 1458 1009 1464
rect 1037 1458 1049 1464
rect 1116 1458 1128 1464
rect 1166 1458 1178 1464
rect 1257 1504 1265 1506
rect 1297 1538 1337 1544
rect 1297 1536 1309 1538
rect 1416 1504 1424 1587
rect 1516 1581 1524 1609
rect 1618 1593 1626 1636
rect 1769 1636 1797 1642
rect 1757 1633 1809 1636
rect 1874 1636 1900 1647
rect 1957 1676 1969 1682
rect 2018 1676 2030 1682
rect 2171 1676 2183 1682
rect 2217 1676 2229 1682
rect 2299 1676 2311 1682
rect 2357 1676 2369 1682
rect 2405 1676 2417 1682
rect 2467 1676 2479 1682
rect 2571 1676 2583 1682
rect 2661 1676 2673 1682
rect 2717 1676 2729 1682
rect 2757 1676 2769 1682
rect 1817 1622 1825 1636
rect 1706 1618 1724 1620
rect 1694 1609 1724 1618
rect 1800 1615 1825 1622
rect 1716 1581 1724 1609
rect 1518 1512 1525 1567
rect 1618 1544 1626 1579
rect 1799 1593 1807 1615
rect 1874 1593 1882 1636
rect 1976 1601 1984 1656
rect 2135 1622 2143 1636
rect 2163 1636 2191 1642
rect 2151 1633 2203 1636
rect 2066 1618 2084 1620
rect 2054 1609 2084 1618
rect 2135 1615 2160 1622
rect 1997 1597 2033 1603
rect 1478 1506 1525 1512
rect 1478 1504 1489 1506
rect 1197 1458 1209 1464
rect 1237 1458 1249 1464
rect 1317 1458 1329 1464
rect 1431 1458 1443 1464
rect 1517 1504 1525 1506
rect 1557 1538 1597 1544
rect 1557 1536 1569 1538
rect 1718 1512 1725 1567
rect 1793 1544 1801 1579
rect 1874 1544 1882 1579
rect 1678 1506 1725 1512
rect 1678 1504 1689 1506
rect 1717 1504 1725 1506
rect 1903 1538 1943 1544
rect 1931 1536 1943 1538
rect 1976 1504 1984 1587
rect 1997 1547 2003 1597
rect 2076 1581 2084 1609
rect 2117 1597 2133 1603
rect 2078 1512 2085 1567
rect 2117 1543 2123 1597
rect 2153 1593 2161 1615
rect 2236 1601 2244 1656
rect 2447 1656 2460 1662
rect 2331 1650 2338 1656
rect 2327 1642 2338 1650
rect 2388 1644 2395 1656
rect 2453 1650 2460 1656
rect 2277 1621 2285 1636
rect 2388 1637 2409 1644
rect 2367 1626 2373 1628
rect 2434 1626 2441 1632
rect 2277 1607 2293 1621
rect 2367 1620 2441 1626
rect 2159 1544 2167 1579
rect 2107 1537 2123 1543
rect 2038 1506 2085 1512
rect 2038 1504 2049 1506
rect 2077 1504 2085 1506
rect 2236 1504 2244 1587
rect 2277 1544 2285 1607
rect 2293 1593 2307 1607
rect 2299 1548 2313 1556
rect 1457 1458 1469 1464
rect 1497 1458 1509 1464
rect 1577 1458 1589 1464
rect 1657 1458 1669 1464
rect 1697 1458 1709 1464
rect 1762 1458 1774 1464
rect 1812 1458 1824 1464
rect 1911 1458 1923 1464
rect 1957 1458 1969 1464
rect 2017 1458 2029 1464
rect 2057 1458 2069 1464
rect 2136 1458 2148 1464
rect 2186 1458 2198 1464
rect 2367 1548 2373 1620
rect 2434 1612 2441 1620
rect 2446 1604 2480 1612
rect 2474 1599 2480 1604
rect 2427 1586 2454 1593
rect 2333 1542 2373 1548
rect 2381 1548 2425 1554
rect 2333 1524 2339 1542
rect 2381 1534 2387 1548
rect 2493 1552 2499 1636
rect 2535 1622 2543 1636
rect 2563 1636 2591 1642
rect 2551 1633 2603 1636
rect 2631 1636 2641 1646
rect 2800 1676 2812 1682
rect 2850 1676 2862 1682
rect 2535 1615 2560 1622
rect 2553 1593 2561 1615
rect 2631 1593 2639 1636
rect 2691 1626 2703 1636
rect 2665 1618 2703 1626
rect 2631 1579 2633 1593
rect 2437 1544 2499 1552
rect 2559 1544 2567 1579
rect 2631 1544 2639 1579
rect 2357 1528 2387 1534
rect 2405 1530 2443 1538
rect 2435 1524 2443 1530
rect 2327 1484 2339 1518
rect 2385 1510 2407 1522
rect 2435 1510 2453 1524
rect 2381 1504 2393 1510
rect 2435 1504 2443 1510
rect 2674 1504 2682 1618
rect 2740 1613 2747 1656
rect 2911 1676 2923 1682
rect 2951 1676 2963 1682
rect 3011 1676 3023 1682
rect 3071 1676 3083 1682
rect 3117 1676 3129 1682
rect 3199 1676 3211 1682
rect 3329 1676 3341 1682
rect 3411 1676 3423 1682
rect 3481 1676 3493 1682
rect 3543 1676 3555 1682
rect 3591 1676 3603 1682
rect 3649 1676 3661 1682
rect 3697 1676 3709 1682
rect 3791 1676 3803 1682
rect 3871 1676 3883 1682
rect 3917 1676 3929 1682
rect 3957 1676 3969 1682
rect 2840 1636 2866 1647
rect 2740 1551 2747 1599
rect 2858 1593 2866 1636
rect 2933 1613 2940 1656
rect 2996 1601 3004 1656
rect 2740 1544 2757 1551
rect 2858 1544 2866 1579
rect 2933 1551 2940 1599
rect 3056 1601 3064 1656
rect 3109 1636 3137 1642
rect 3097 1633 3149 1636
rect 3157 1622 3165 1636
rect 3229 1628 3241 1636
rect 3140 1615 3165 1622
rect 3217 1622 3241 1628
rect 3299 1628 3311 1636
rect 3299 1622 3323 1628
rect 2923 1544 2940 1551
rect 2217 1458 2229 1464
rect 2297 1458 2309 1464
rect 2355 1458 2367 1464
rect 2401 1458 2413 1464
rect 2467 1458 2479 1464
rect 2536 1458 2548 1464
rect 2586 1458 2598 1464
rect 2647 1458 2659 1464
rect 2691 1458 2703 1464
rect 2797 1538 2837 1544
rect 2797 1536 2809 1538
rect 2996 1504 3004 1587
rect 3056 1504 3064 1587
rect 3139 1593 3147 1615
rect 3133 1544 3141 1579
rect 3217 1573 3225 1622
rect 3315 1573 3323 1622
rect 3375 1622 3383 1636
rect 3403 1636 3431 1642
rect 3391 1633 3443 1636
rect 3500 1656 3513 1662
rect 3500 1650 3507 1656
rect 3565 1644 3572 1656
rect 3375 1615 3400 1622
rect 3357 1597 3373 1603
rect 2717 1458 2729 1464
rect 2817 1458 2829 1464
rect 2951 1458 2963 1464
rect 3011 1458 3023 1464
rect 3071 1458 3083 1464
rect 3217 1504 3225 1559
rect 3315 1504 3323 1559
rect 3357 1523 3363 1597
rect 3393 1593 3401 1615
rect 3399 1544 3407 1579
rect 3461 1552 3467 1636
rect 3551 1637 3572 1644
rect 3622 1650 3629 1656
rect 3622 1642 3633 1650
rect 3519 1626 3526 1632
rect 3587 1626 3593 1628
rect 3519 1620 3593 1626
rect 3675 1621 3683 1636
rect 3519 1612 3526 1620
rect 3480 1604 3514 1612
rect 3480 1599 3486 1604
rect 3506 1586 3533 1593
rect 3461 1544 3523 1552
rect 3535 1548 3579 1554
rect 3357 1517 3373 1523
rect 3102 1458 3114 1464
rect 3152 1458 3164 1464
rect 3197 1458 3209 1464
rect 3237 1458 3249 1464
rect 3291 1458 3303 1464
rect 3331 1458 3343 1464
rect 3517 1530 3555 1538
rect 3573 1534 3579 1548
rect 3587 1548 3593 1620
rect 3667 1607 3683 1621
rect 3653 1593 3667 1607
rect 3587 1542 3627 1548
rect 3647 1548 3661 1556
rect 3675 1544 3683 1607
rect 3716 1601 3724 1656
rect 3776 1601 3784 1656
rect 3835 1622 3843 1636
rect 3863 1636 3891 1642
rect 3997 1676 4009 1682
rect 4037 1676 4049 1682
rect 4077 1676 4089 1682
rect 4140 1676 4152 1682
rect 4190 1676 4202 1682
rect 3851 1633 3903 1636
rect 3835 1615 3860 1622
rect 3853 1593 3861 1615
rect 3940 1613 3947 1656
rect 4020 1613 4027 1656
rect 3517 1524 3525 1530
rect 3573 1528 3603 1534
rect 3621 1524 3627 1542
rect 3507 1510 3525 1524
rect 3553 1510 3575 1522
rect 3517 1504 3525 1510
rect 3567 1504 3579 1510
rect 3621 1484 3633 1518
rect 3716 1504 3724 1587
rect 3776 1504 3784 1587
rect 4096 1601 4104 1656
rect 4237 1676 4249 1682
rect 4277 1676 4289 1682
rect 4320 1676 4332 1682
rect 4370 1676 4382 1682
rect 4180 1636 4206 1647
rect 3859 1544 3867 1579
rect 3940 1551 3947 1599
rect 4020 1551 4027 1599
rect 4198 1593 4206 1636
rect 4260 1613 4267 1656
rect 4417 1676 4429 1682
rect 4477 1676 4489 1682
rect 4571 1676 4583 1682
rect 4617 1676 4629 1682
rect 4699 1676 4711 1682
rect 4360 1636 4386 1647
rect 3940 1544 3957 1551
rect 4020 1544 4037 1551
rect 3376 1458 3388 1464
rect 3426 1458 3438 1464
rect 3481 1458 3493 1464
rect 3547 1458 3559 1464
rect 3593 1458 3605 1464
rect 3651 1458 3663 1464
rect 3697 1458 3709 1464
rect 3791 1458 3803 1464
rect 3836 1458 3848 1464
rect 3886 1458 3898 1464
rect 4096 1504 4104 1587
rect 4198 1544 4206 1579
rect 4217 1567 4223 1613
rect 4260 1551 4267 1599
rect 4378 1593 4386 1636
rect 4436 1601 4444 1656
rect 4496 1601 4504 1656
rect 4556 1601 4564 1656
rect 4609 1636 4637 1642
rect 4597 1633 4649 1636
rect 4657 1622 4665 1636
rect 4729 1628 4741 1636
rect 4640 1615 4665 1622
rect 4260 1544 4277 1551
rect 4378 1544 4386 1579
rect 4137 1538 4177 1544
rect 4137 1536 4149 1538
rect 4317 1538 4357 1544
rect 4317 1536 4329 1538
rect 4436 1504 4444 1587
rect 4496 1504 4504 1587
rect 4556 1504 4564 1587
rect 4639 1593 4647 1615
rect 4717 1622 4741 1628
rect 4633 1544 4641 1579
rect 3917 1458 3929 1464
rect 3997 1458 4009 1464
rect 4077 1458 4089 1464
rect 4157 1458 4169 1464
rect 4237 1458 4249 1464
rect 4337 1458 4349 1464
rect 4417 1458 4429 1464
rect 4477 1458 4489 1464
rect 4571 1458 4583 1464
rect 4677 1523 4683 1613
rect 4717 1573 4725 1622
rect 4667 1517 4683 1523
rect 4717 1504 4725 1559
rect 4602 1458 4614 1464
rect 4652 1458 4664 1464
rect 4697 1458 4709 1464
rect 4737 1458 4749 1464
rect -62 1456 4776 1458
rect -62 1444 4 1456
rect -62 1442 4776 1444
rect -62 978 -2 1442
rect 71 1436 83 1442
rect 117 1436 129 1442
rect 157 1436 169 1442
rect 217 1436 229 1442
rect 257 1436 269 1442
rect 331 1436 343 1442
rect 371 1436 383 1442
rect 138 1394 149 1396
rect 177 1394 185 1396
rect 138 1388 185 1394
rect 238 1394 249 1396
rect 402 1436 414 1442
rect 452 1436 464 1442
rect 517 1436 529 1442
rect 602 1436 614 1442
rect 652 1436 664 1442
rect 277 1394 285 1396
rect 238 1388 285 1394
rect 91 1362 103 1364
rect 63 1356 103 1362
rect 34 1321 42 1356
rect 178 1333 185 1388
rect 34 1264 42 1307
rect 176 1291 184 1319
rect 197 1303 203 1353
rect 278 1333 285 1388
rect 197 1297 213 1303
rect 276 1291 284 1319
rect 34 1253 60 1264
rect 38 1218 50 1224
rect 88 1218 100 1224
rect 154 1282 184 1291
rect 166 1280 184 1282
rect 254 1282 284 1291
rect 297 1287 303 1353
rect 355 1341 363 1396
rect 266 1280 284 1282
rect 355 1278 363 1327
rect 433 1321 441 1356
rect 497 1362 509 1364
rect 497 1356 537 1362
rect 702 1436 714 1442
rect 752 1436 764 1442
rect 797 1436 809 1442
rect 841 1436 853 1442
rect 911 1436 923 1442
rect 951 1436 963 1442
rect 477 1307 483 1353
rect 558 1321 566 1356
rect 633 1321 641 1356
rect 733 1321 741 1356
rect 439 1285 447 1307
rect 440 1278 465 1285
rect 339 1272 363 1278
rect 339 1264 351 1272
rect 397 1264 449 1267
rect 409 1258 437 1264
rect 457 1264 465 1278
rect 558 1264 566 1307
rect 639 1285 647 1307
rect 739 1285 747 1307
rect 640 1278 665 1285
rect 740 1278 765 1285
rect 818 1282 826 1396
rect 977 1436 989 1442
rect 1017 1436 1029 1442
rect 1091 1436 1103 1442
rect 1131 1436 1143 1442
rect 1191 1436 1203 1442
rect 1247 1436 1259 1442
rect 1291 1436 1303 1442
rect 861 1321 869 1356
rect 935 1341 943 1396
rect 997 1341 1005 1396
rect 1075 1394 1083 1396
rect 1111 1394 1122 1396
rect 1075 1388 1122 1394
rect 867 1307 869 1321
rect 540 1253 566 1264
rect 597 1264 649 1267
rect 609 1258 637 1264
rect 657 1264 665 1278
rect 697 1264 749 1267
rect 709 1258 737 1264
rect 757 1264 765 1278
rect 797 1274 835 1282
rect 797 1264 809 1274
rect 861 1264 869 1307
rect 935 1278 943 1327
rect 1075 1333 1082 1388
rect 859 1254 869 1264
rect 919 1272 943 1278
rect 997 1278 1005 1327
rect 1076 1291 1084 1319
rect 1176 1313 1184 1396
rect 1322 1436 1334 1442
rect 1372 1436 1384 1442
rect 1231 1321 1239 1356
rect 1231 1307 1233 1321
rect 1076 1282 1106 1291
rect 1076 1280 1094 1282
rect 997 1272 1021 1278
rect 919 1264 931 1272
rect 1009 1264 1021 1272
rect 118 1218 130 1224
rect 218 1218 230 1224
rect 369 1218 381 1224
rect 417 1218 429 1224
rect 500 1218 512 1224
rect 550 1218 562 1224
rect 617 1218 629 1224
rect 717 1218 729 1224
rect 827 1218 839 1224
rect 949 1218 961 1224
rect 1176 1244 1184 1299
rect 1231 1264 1239 1307
rect 1274 1282 1282 1396
rect 1436 1436 1448 1442
rect 1486 1436 1498 1442
rect 1417 1377 1433 1383
rect 1353 1321 1361 1356
rect 1359 1285 1367 1307
rect 1417 1303 1423 1377
rect 1517 1436 1529 1442
rect 1557 1436 1569 1442
rect 1602 1436 1614 1442
rect 1652 1436 1664 1442
rect 1459 1321 1467 1356
rect 1537 1341 1545 1396
rect 1697 1436 1709 1442
rect 1737 1436 1749 1442
rect 1797 1436 1809 1442
rect 1877 1436 1889 1442
rect 1917 1436 1929 1442
rect 1982 1436 1994 1442
rect 2032 1436 2044 1442
rect 1417 1297 1433 1303
rect 1453 1285 1461 1307
rect 1265 1274 1303 1282
rect 1360 1278 1385 1285
rect 1291 1264 1303 1274
rect 1231 1254 1241 1264
rect 1317 1264 1369 1267
rect 1329 1258 1357 1264
rect 1377 1264 1385 1278
rect 1435 1278 1460 1285
rect 1537 1278 1545 1327
rect 1633 1321 1641 1356
rect 1717 1341 1725 1396
rect 1777 1362 1789 1364
rect 1777 1356 1817 1362
rect 1898 1394 1909 1396
rect 1937 1394 1945 1396
rect 1898 1388 1945 1394
rect 1639 1285 1647 1307
rect 1640 1278 1665 1285
rect 1435 1264 1443 1278
rect 1537 1272 1561 1278
rect 1451 1264 1503 1267
rect 1549 1264 1561 1272
rect 1463 1258 1491 1264
rect 1597 1264 1649 1267
rect 1609 1258 1637 1264
rect 1657 1264 1665 1278
rect 1717 1278 1725 1327
rect 1838 1321 1846 1356
rect 1938 1333 1945 1388
rect 2077 1436 2089 1442
rect 2137 1436 2149 1442
rect 2177 1436 2189 1442
rect 2237 1436 2249 1442
rect 2277 1436 2289 1442
rect 2347 1436 2359 1442
rect 2431 1436 2443 1442
rect 2471 1436 2483 1442
rect 2013 1321 2021 1356
rect 1717 1272 1741 1278
rect 1729 1264 1741 1272
rect 1838 1264 1846 1307
rect 1936 1291 1944 1319
rect 2096 1313 2104 1396
rect 2158 1394 2169 1396
rect 2197 1394 2205 1396
rect 2158 1388 2205 1394
rect 2198 1333 2205 1388
rect 2257 1341 2265 1396
rect 2497 1436 2509 1442
rect 2589 1436 2601 1442
rect 2642 1436 2654 1442
rect 2692 1436 2704 1442
rect 2379 1357 2383 1366
rect 2317 1348 2325 1356
rect 2317 1340 2353 1348
rect 1820 1253 1846 1264
rect 979 1218 991 1224
rect 1130 1218 1142 1224
rect 1191 1218 1203 1224
rect 1261 1218 1273 1224
rect 1337 1218 1349 1224
rect 1471 1218 1483 1224
rect 1519 1218 1531 1224
rect 1617 1218 1629 1224
rect 1699 1218 1711 1224
rect 1780 1218 1792 1224
rect 1830 1218 1842 1224
rect 1914 1282 1944 1291
rect 2019 1285 2027 1307
rect 1926 1280 1944 1282
rect 2020 1278 2045 1285
rect 1977 1264 2029 1267
rect 1989 1258 2017 1264
rect 2037 1264 2045 1278
rect 2096 1244 2104 1299
rect 2196 1291 2204 1319
rect 2174 1282 2204 1291
rect 2186 1280 2204 1282
rect 2257 1278 2265 1327
rect 2358 1284 2364 1339
rect 2374 1313 2383 1357
rect 2455 1341 2463 1396
rect 2257 1272 2281 1278
rect 2269 1264 2281 1272
rect 2343 1272 2353 1278
rect 2343 1244 2349 1272
rect 2380 1264 2387 1299
rect 2455 1278 2463 1327
rect 2516 1313 2524 1396
rect 2571 1321 2579 1356
rect 2615 1350 2623 1396
rect 2761 1436 2773 1442
rect 2831 1436 2843 1442
rect 2881 1436 2893 1442
rect 2947 1436 2959 1442
rect 2993 1436 3005 1442
rect 3051 1436 3063 1442
rect 3151 1436 3163 1442
rect 3231 1436 3243 1442
rect 3301 1436 3313 1442
rect 3367 1436 3379 1442
rect 3413 1436 3425 1442
rect 3471 1436 3483 1442
rect 3551 1436 3563 1442
rect 3631 1436 3643 1442
rect 3711 1436 3723 1442
rect 2917 1390 2925 1396
rect 2967 1390 2979 1396
rect 2907 1376 2925 1390
rect 2953 1378 2975 1390
rect 3021 1382 3033 1416
rect 2917 1370 2925 1376
rect 2917 1362 2955 1370
rect 2973 1366 3003 1372
rect 2597 1344 2623 1350
rect 2597 1338 2600 1344
rect 2571 1307 2573 1321
rect 2439 1272 2463 1278
rect 2439 1264 2451 1272
rect 2516 1244 2524 1299
rect 2571 1264 2579 1307
rect 2593 1282 2600 1338
rect 2673 1321 2681 1356
rect 2795 1321 2803 1356
rect 2861 1348 2923 1356
rect 2679 1285 2687 1307
rect 2597 1276 2600 1282
rect 2680 1278 2705 1285
rect 2796 1281 2804 1307
rect 2597 1270 2619 1276
rect 1878 1218 1890 1224
rect 1997 1218 2009 1224
rect 2077 1218 2089 1224
rect 2138 1218 2150 1224
rect 2239 1218 2251 1224
rect 2317 1218 2325 1224
rect 2357 1218 2369 1224
rect 2469 1218 2481 1224
rect 2611 1244 2619 1270
rect 2637 1264 2689 1267
rect 2649 1258 2677 1264
rect 2697 1264 2705 1278
rect 2775 1274 2804 1281
rect 2775 1264 2781 1274
rect 2791 1264 2843 1266
rect 2763 1224 2791 1230
rect 2803 1260 2831 1264
rect 2861 1264 2867 1348
rect 2973 1352 2979 1366
rect 3021 1358 3027 1376
rect 2935 1346 2979 1352
rect 2987 1352 3027 1358
rect 2906 1307 2933 1314
rect 2880 1296 2886 1301
rect 2880 1288 2914 1296
rect 2919 1280 2926 1288
rect 2987 1280 2993 1352
rect 3047 1344 3061 1352
rect 3053 1293 3067 1307
rect 3075 1293 3083 1356
rect 3251 1362 3263 1364
rect 3223 1356 3263 1362
rect 3337 1390 3345 1396
rect 3387 1390 3399 1396
rect 3327 1376 3345 1390
rect 3373 1378 3395 1390
rect 3441 1382 3453 1416
rect 3337 1370 3345 1376
rect 3337 1362 3375 1370
rect 3393 1366 3423 1372
rect 3123 1349 3140 1356
rect 2919 1274 2993 1280
rect 3067 1279 3083 1293
rect 2919 1268 2926 1274
rect 2987 1272 2993 1274
rect 2951 1256 2972 1263
rect 3075 1264 3083 1279
rect 2900 1244 2907 1250
rect 2965 1244 2972 1256
rect 3022 1250 3033 1258
rect 3022 1244 3029 1250
rect 2900 1238 2913 1244
rect 3133 1301 3140 1349
rect 3194 1321 3202 1356
rect 3281 1348 3343 1356
rect 3133 1244 3140 1287
rect 3194 1264 3202 1307
rect 3281 1264 3287 1348
rect 3393 1352 3399 1366
rect 3441 1358 3447 1376
rect 3355 1346 3399 1352
rect 3407 1352 3447 1358
rect 3326 1307 3353 1314
rect 3300 1296 3306 1301
rect 3300 1288 3334 1296
rect 3339 1280 3346 1288
rect 3407 1280 3413 1352
rect 3467 1344 3481 1352
rect 3473 1293 3487 1307
rect 3495 1293 3503 1356
rect 3536 1313 3544 1396
rect 3737 1436 3749 1442
rect 3817 1436 3829 1442
rect 3875 1436 3887 1442
rect 3921 1436 3933 1442
rect 3987 1436 3999 1442
rect 4042 1436 4054 1442
rect 4092 1436 4104 1442
rect 3603 1349 3620 1356
rect 3683 1349 3700 1356
rect 3613 1301 3620 1349
rect 3693 1301 3700 1349
rect 3756 1313 3764 1396
rect 3847 1382 3859 1416
rect 3901 1390 3913 1396
rect 3955 1390 3963 1396
rect 3905 1378 3927 1390
rect 3955 1376 3973 1390
rect 3853 1358 3859 1376
rect 3877 1366 3907 1372
rect 3955 1370 3963 1376
rect 3339 1274 3413 1280
rect 3487 1279 3503 1293
rect 3339 1268 3346 1274
rect 3407 1272 3413 1274
rect 3194 1253 3220 1264
rect 2497 1218 2509 1224
rect 2589 1218 2601 1224
rect 2657 1218 2669 1224
rect 2811 1218 2823 1224
rect 2881 1218 2893 1224
rect 2943 1218 2955 1224
rect 2991 1218 3003 1224
rect 3049 1218 3061 1224
rect 3111 1218 3123 1224
rect 3151 1218 3163 1224
rect 3371 1256 3392 1263
rect 3495 1264 3503 1279
rect 3320 1244 3327 1250
rect 3385 1244 3392 1256
rect 3442 1250 3453 1258
rect 3442 1244 3449 1250
rect 3320 1238 3333 1244
rect 3536 1244 3544 1299
rect 3613 1244 3620 1287
rect 3693 1244 3700 1287
rect 3756 1244 3764 1299
rect 3797 1293 3805 1356
rect 3819 1344 3833 1352
rect 3853 1352 3893 1358
rect 3813 1293 3827 1307
rect 3797 1279 3813 1293
rect 3887 1280 3893 1352
rect 3901 1352 3907 1366
rect 3925 1362 3963 1370
rect 4137 1436 4149 1442
rect 4177 1436 4189 1442
rect 4249 1436 4261 1442
rect 4311 1436 4323 1442
rect 4351 1436 4363 1442
rect 3901 1346 3945 1352
rect 3957 1348 4019 1356
rect 3947 1307 3974 1314
rect 3994 1296 4000 1301
rect 3966 1288 4000 1296
rect 3954 1280 3961 1288
rect 3797 1264 3805 1279
rect 3887 1274 3961 1280
rect 3887 1272 3893 1274
rect 3198 1218 3210 1224
rect 3248 1218 3260 1224
rect 3301 1218 3313 1224
rect 3363 1218 3375 1224
rect 3411 1218 3423 1224
rect 3469 1218 3481 1224
rect 3551 1218 3563 1224
rect 3591 1218 3603 1224
rect 3631 1218 3643 1224
rect 3671 1218 3683 1224
rect 3711 1218 3723 1224
rect 3954 1268 3961 1274
rect 3847 1250 3858 1258
rect 3851 1244 3858 1250
rect 3908 1256 3929 1263
rect 4013 1264 4019 1348
rect 4073 1321 4081 1356
rect 4157 1341 4165 1396
rect 4396 1436 4408 1442
rect 4446 1436 4458 1442
rect 4079 1285 4087 1307
rect 4080 1278 4105 1285
rect 3908 1244 3915 1256
rect 3973 1244 3980 1250
rect 3967 1238 3980 1244
rect 4037 1264 4089 1267
rect 4049 1258 4077 1264
rect 4097 1264 4105 1278
rect 4157 1278 4165 1327
rect 4231 1321 4239 1356
rect 4275 1350 4283 1396
rect 4257 1344 4283 1350
rect 4257 1338 4260 1344
rect 4335 1341 4343 1396
rect 4496 1436 4508 1442
rect 4546 1436 4558 1442
rect 4577 1436 4589 1442
rect 4657 1436 4669 1442
rect 4751 1436 4763 1442
rect 4231 1307 4233 1321
rect 4157 1272 4181 1278
rect 4169 1264 4181 1272
rect 4231 1264 4239 1307
rect 4253 1282 4260 1338
rect 4257 1276 4260 1282
rect 4335 1278 4343 1327
rect 4419 1321 4427 1356
rect 4519 1321 4527 1356
rect 4600 1349 4617 1356
rect 4413 1285 4421 1307
rect 4513 1285 4521 1307
rect 4600 1301 4607 1349
rect 4676 1313 4684 1396
rect 4736 1313 4744 1396
rect 4257 1270 4279 1276
rect 4271 1244 4279 1270
rect 4319 1272 4343 1278
rect 4395 1278 4420 1285
rect 4495 1278 4520 1285
rect 4319 1264 4331 1272
rect 4395 1264 4403 1278
rect 4411 1264 4463 1267
rect 4495 1264 4503 1278
rect 4423 1258 4451 1264
rect 4511 1264 4563 1267
rect 4523 1258 4551 1264
rect 4600 1244 4607 1287
rect 4676 1244 4684 1299
rect 4736 1244 4744 1299
rect 3737 1218 3749 1224
rect 3819 1218 3831 1224
rect 3877 1218 3889 1224
rect 3925 1218 3937 1224
rect 3987 1218 3999 1224
rect 4057 1218 4069 1224
rect 4139 1218 4151 1224
rect 4249 1218 4261 1224
rect 4349 1218 4361 1224
rect 4431 1218 4443 1224
rect 4531 1218 4543 1224
rect 4577 1218 4589 1224
rect 4617 1218 4629 1224
rect 4657 1218 4669 1224
rect 4751 1218 4763 1224
rect 4782 1218 4842 1682
rect 4 1216 4842 1218
rect 4776 1204 4842 1216
rect 4 1202 4842 1204
rect 71 1196 83 1202
rect 137 1196 149 1202
rect 218 1196 230 1202
rect 320 1196 332 1202
rect 370 1196 382 1202
rect 35 1142 43 1156
rect 63 1156 91 1162
rect 51 1153 103 1156
rect 129 1156 157 1162
rect 117 1153 169 1156
rect 177 1142 185 1156
rect 35 1135 60 1142
rect 160 1135 185 1142
rect 418 1196 430 1202
rect 520 1196 532 1202
rect 570 1196 582 1202
rect 669 1196 681 1202
rect 741 1196 753 1202
rect 870 1196 882 1202
rect 951 1196 963 1202
rect 1017 1196 1029 1202
rect 1151 1196 1163 1202
rect 1249 1196 1261 1202
rect 1321 1196 1333 1202
rect 1379 1196 1391 1202
rect 1491 1196 1503 1202
rect 1569 1196 1581 1202
rect 1649 1196 1661 1202
rect 360 1156 386 1167
rect 266 1138 284 1140
rect 53 1113 61 1135
rect 159 1113 167 1135
rect 254 1129 284 1138
rect 276 1101 284 1129
rect 59 1064 67 1099
rect 153 1064 161 1099
rect 297 1087 303 1133
rect 378 1113 386 1156
rect 487 1157 503 1163
rect 466 1138 484 1140
rect 454 1129 484 1138
rect 476 1101 484 1129
rect 36 978 48 984
rect 86 978 98 984
rect 278 1032 285 1087
rect 378 1064 386 1099
rect 238 1026 285 1032
rect 238 1024 249 1026
rect 122 978 134 984
rect 172 978 184 984
rect 277 1024 285 1026
rect 317 1058 357 1064
rect 317 1056 329 1058
rect 478 1032 485 1087
rect 497 1083 503 1157
rect 560 1156 586 1167
rect 578 1113 586 1156
rect 711 1156 721 1166
rect 639 1148 651 1156
rect 639 1142 663 1148
rect 497 1077 513 1083
rect 578 1064 586 1099
rect 655 1093 663 1142
rect 711 1113 719 1156
rect 771 1146 783 1156
rect 745 1138 783 1146
rect 816 1138 834 1140
rect 711 1099 713 1113
rect 438 1026 485 1032
rect 438 1024 449 1026
rect 477 1024 485 1026
rect 517 1058 557 1064
rect 517 1056 529 1058
rect 655 1024 663 1079
rect 711 1064 719 1099
rect 754 1024 762 1138
rect 816 1129 846 1138
rect 915 1142 923 1156
rect 943 1156 971 1162
rect 931 1153 983 1156
rect 1009 1156 1037 1162
rect 997 1153 1049 1156
rect 1057 1142 1065 1156
rect 915 1135 940 1142
rect 1040 1135 1065 1142
rect 1115 1142 1123 1156
rect 1143 1156 1171 1162
rect 1131 1153 1183 1156
rect 1291 1156 1301 1166
rect 1678 1196 1690 1202
rect 1829 1196 1841 1202
rect 1219 1148 1231 1156
rect 1219 1142 1243 1148
rect 1115 1135 1140 1142
rect 816 1101 824 1129
rect 867 1117 903 1123
rect 815 1032 822 1087
rect 897 1047 903 1117
rect 933 1113 941 1135
rect 1039 1113 1047 1135
rect 1133 1113 1141 1135
rect 939 1064 947 1099
rect 1033 1064 1041 1099
rect 1139 1064 1147 1099
rect 1235 1093 1243 1142
rect 1291 1113 1299 1156
rect 1351 1146 1363 1156
rect 1409 1148 1421 1156
rect 1325 1138 1363 1146
rect 1397 1142 1421 1148
rect 1291 1099 1293 1113
rect 815 1026 862 1032
rect 815 1024 823 1026
rect 851 1024 862 1026
rect 217 978 229 984
rect 257 978 269 984
rect 337 978 349 984
rect 417 978 429 984
rect 457 978 469 984
rect 537 978 549 984
rect 631 978 643 984
rect 671 978 683 984
rect 727 978 739 984
rect 771 978 783 984
rect 831 978 843 984
rect 871 978 883 984
rect 916 978 928 984
rect 966 978 978 984
rect 1002 978 1014 984
rect 1052 978 1064 984
rect 1235 1024 1243 1079
rect 1291 1064 1299 1099
rect 1116 978 1128 984
rect 1166 978 1178 984
rect 1334 1024 1342 1138
rect 1397 1093 1405 1142
rect 1476 1113 1484 1156
rect 1539 1148 1551 1156
rect 1619 1148 1631 1156
rect 1539 1142 1563 1148
rect 1397 1024 1405 1079
rect 1476 1064 1484 1099
rect 1555 1093 1563 1142
rect 1587 1137 1603 1143
rect 1619 1142 1643 1148
rect 1211 978 1223 984
rect 1251 978 1263 984
rect 1307 978 1319 984
rect 1351 978 1363 984
rect 1555 1024 1563 1079
rect 1597 1063 1603 1137
rect 1635 1093 1643 1142
rect 1858 1196 1870 1202
rect 1959 1196 1971 1202
rect 2072 1196 2084 1202
rect 2128 1196 2140 1202
rect 2230 1196 2242 1202
rect 2309 1196 2321 1202
rect 1799 1148 1811 1156
rect 1799 1142 1823 1148
rect 1726 1138 1744 1140
rect 1714 1129 1744 1138
rect 1736 1101 1744 1129
rect 1815 1093 1823 1142
rect 1989 1148 2001 1156
rect 1977 1142 2001 1148
rect 1906 1138 1924 1140
rect 1894 1129 1924 1138
rect 1916 1101 1924 1129
rect 1597 1057 1623 1063
rect 1617 1047 1623 1057
rect 1635 1024 1643 1079
rect 1738 1032 1745 1087
rect 1977 1093 1985 1142
rect 1698 1026 1745 1032
rect 1698 1024 1709 1026
rect 1377 978 1389 984
rect 1417 978 1429 984
rect 1491 978 1503 984
rect 1531 978 1543 984
rect 1571 978 1583 984
rect 1611 978 1623 984
rect 1651 978 1663 984
rect 1737 1024 1745 1026
rect 1815 1024 1823 1079
rect 1918 1032 1925 1087
rect 2100 1113 2107 1156
rect 2176 1138 2194 1140
rect 2176 1129 2206 1138
rect 2340 1196 2352 1202
rect 2390 1196 2402 1202
rect 2471 1196 2483 1202
rect 2549 1196 2561 1202
rect 2651 1196 2663 1202
rect 2719 1196 2731 1202
rect 2801 1196 2813 1202
rect 2863 1196 2875 1202
rect 2911 1196 2923 1202
rect 2969 1196 2981 1202
rect 3019 1196 3031 1202
rect 3151 1196 3163 1202
rect 3197 1196 3209 1202
rect 3237 1196 3249 1202
rect 3277 1196 3289 1202
rect 3349 1196 3361 1202
rect 3419 1196 3431 1202
rect 3477 1196 3489 1202
rect 3517 1196 3529 1202
rect 3557 1196 3569 1202
rect 3597 1196 3609 1202
rect 3637 1196 3649 1202
rect 2380 1156 2406 1167
rect 2279 1148 2291 1156
rect 2279 1142 2303 1148
rect 2176 1101 2184 1129
rect 2227 1117 2263 1123
rect 1878 1026 1925 1032
rect 1878 1024 1889 1026
rect 1677 978 1689 984
rect 1717 978 1729 984
rect 1791 978 1803 984
rect 1831 978 1843 984
rect 1917 1024 1925 1026
rect 1977 1024 1985 1079
rect 2093 1076 2099 1099
rect 2072 1070 2099 1076
rect 2072 1064 2084 1070
rect 2063 984 2091 990
rect 2103 1056 2131 1062
rect 2175 1032 2182 1087
rect 2257 1063 2263 1117
rect 2295 1093 2303 1142
rect 2398 1113 2406 1156
rect 2456 1121 2464 1176
rect 2603 1190 2631 1196
rect 2643 1156 2671 1160
rect 2519 1148 2531 1156
rect 2519 1142 2543 1148
rect 2257 1057 2273 1063
rect 2175 1026 2222 1032
rect 2175 1024 2183 1026
rect 2211 1024 2222 1026
rect 2295 1024 2303 1079
rect 2398 1064 2406 1099
rect 2337 1058 2377 1064
rect 2337 1056 2349 1058
rect 1857 978 1869 984
rect 1897 978 1909 984
rect 1957 978 1969 984
rect 1997 978 2009 984
rect 2111 978 2123 984
rect 2191 978 2203 984
rect 2231 978 2243 984
rect 2456 1024 2464 1107
rect 2535 1093 2543 1142
rect 2615 1146 2621 1156
rect 2631 1154 2683 1156
rect 2701 1150 2709 1176
rect 2820 1176 2833 1182
rect 2820 1170 2827 1176
rect 2885 1164 2892 1176
rect 2615 1139 2644 1146
rect 2701 1144 2723 1150
rect 2636 1113 2644 1139
rect 2720 1138 2723 1144
rect 2535 1024 2543 1079
rect 2635 1064 2643 1099
rect 2720 1082 2727 1138
rect 2741 1113 2749 1156
rect 2747 1099 2749 1113
rect 2720 1076 2723 1082
rect 2697 1070 2723 1076
rect 2271 978 2283 984
rect 2311 978 2323 984
rect 2357 978 2369 984
rect 2471 978 2483 984
rect 2511 978 2523 984
rect 2551 978 2563 984
rect 2697 1024 2705 1070
rect 2741 1064 2749 1099
rect 2781 1072 2787 1156
rect 2871 1157 2892 1164
rect 2942 1170 2949 1176
rect 2942 1162 2953 1170
rect 2839 1146 2846 1152
rect 2907 1146 2913 1148
rect 2839 1140 2913 1146
rect 2995 1141 3003 1156
rect 3049 1148 3061 1156
rect 2839 1132 2846 1140
rect 2800 1124 2834 1132
rect 2800 1119 2806 1124
rect 2826 1106 2853 1113
rect 2781 1064 2843 1072
rect 2855 1068 2899 1074
rect 2837 1050 2875 1058
rect 2893 1054 2899 1068
rect 2907 1068 2913 1140
rect 2987 1127 3003 1141
rect 2973 1113 2987 1127
rect 2907 1062 2947 1068
rect 2967 1068 2981 1076
rect 2995 1064 3003 1127
rect 3037 1142 3061 1148
rect 3115 1142 3123 1156
rect 3143 1156 3171 1162
rect 3131 1153 3183 1156
rect 3217 1150 3225 1156
rect 3257 1150 3265 1156
rect 3217 1142 3265 1150
rect 3037 1093 3045 1142
rect 3115 1135 3140 1142
rect 3133 1113 3141 1135
rect 3257 1113 3265 1142
rect 3331 1113 3339 1156
rect 3371 1150 3379 1176
rect 3357 1144 3379 1150
rect 3401 1150 3409 1176
rect 3677 1196 3689 1202
rect 3717 1196 3729 1202
rect 3757 1196 3769 1202
rect 3797 1196 3809 1202
rect 3837 1196 3849 1202
rect 3899 1196 3911 1202
rect 3959 1196 3971 1202
rect 4059 1196 4071 1202
rect 4117 1196 4129 1202
rect 4165 1196 4177 1202
rect 4227 1196 4239 1202
rect 4279 1196 4291 1202
rect 4377 1196 4389 1202
rect 4509 1196 4521 1202
rect 4557 1196 4569 1202
rect 4638 1196 4650 1202
rect 3401 1144 3423 1150
rect 3357 1138 3360 1144
rect 3331 1099 3333 1113
rect 2837 1044 2845 1050
rect 2893 1048 2923 1054
rect 2941 1044 2947 1062
rect 2827 1030 2845 1044
rect 2873 1030 2895 1042
rect 2837 1024 2845 1030
rect 2887 1024 2899 1030
rect 2941 1004 2953 1038
rect 3037 1024 3045 1079
rect 3139 1064 3147 1099
rect 3257 1076 3265 1099
rect 3217 1070 3265 1076
rect 3217 1064 3229 1070
rect 3257 1064 3265 1070
rect 3331 1064 3339 1099
rect 3353 1082 3360 1138
rect 3420 1138 3423 1144
rect 3357 1076 3360 1082
rect 3420 1082 3427 1138
rect 3441 1113 3449 1156
rect 3496 1150 3508 1156
rect 3537 1150 3549 1156
rect 3576 1150 3588 1156
rect 3616 1150 3628 1156
rect 3696 1150 3708 1156
rect 3737 1150 3749 1156
rect 3776 1150 3788 1156
rect 3816 1150 3828 1156
rect 3881 1150 3889 1176
rect 3496 1142 3523 1150
rect 3537 1142 3562 1150
rect 3576 1142 3602 1150
rect 3616 1149 3634 1150
rect 3616 1142 3635 1149
rect 3696 1142 3723 1150
rect 3737 1142 3762 1150
rect 3776 1142 3802 1150
rect 3816 1149 3834 1150
rect 3816 1142 3835 1149
rect 3881 1144 3903 1150
rect 3515 1136 3523 1142
rect 3554 1136 3562 1142
rect 3594 1136 3602 1142
rect 3515 1124 3530 1136
rect 3554 1124 3570 1136
rect 3594 1124 3610 1136
rect 3447 1099 3449 1113
rect 3420 1076 3423 1082
rect 3357 1070 3383 1076
rect 2601 978 2613 984
rect 2671 978 2683 984
rect 2719 978 2731 984
rect 2801 978 2813 984
rect 2867 978 2879 984
rect 2913 978 2925 984
rect 2971 978 2983 984
rect 3017 978 3029 984
rect 3057 978 3069 984
rect 3116 978 3128 984
rect 3166 978 3178 984
rect 3375 1024 3383 1070
rect 3397 1070 3423 1076
rect 3397 1024 3405 1070
rect 3441 1064 3449 1099
rect 3515 1078 3523 1124
rect 3554 1078 3562 1124
rect 3594 1078 3602 1124
rect 3628 1121 3635 1142
rect 3715 1136 3723 1142
rect 3754 1136 3762 1142
rect 3794 1136 3802 1142
rect 3715 1124 3730 1136
rect 3754 1124 3770 1136
rect 3794 1124 3810 1136
rect 3628 1107 3633 1121
rect 3628 1078 3635 1107
rect 3715 1078 3723 1124
rect 3754 1078 3762 1124
rect 3794 1078 3802 1124
rect 3828 1121 3835 1142
rect 3900 1138 3903 1144
rect 3828 1107 3833 1121
rect 3828 1078 3835 1107
rect 3497 1070 3523 1078
rect 3537 1070 3562 1078
rect 3577 1070 3602 1078
rect 3617 1070 3635 1078
rect 3697 1070 3723 1078
rect 3737 1070 3762 1078
rect 3777 1070 3802 1078
rect 3817 1070 3835 1078
rect 3900 1082 3907 1138
rect 3921 1113 3929 1156
rect 3989 1148 4001 1156
rect 3977 1142 4001 1148
rect 4207 1176 4220 1182
rect 4091 1170 4098 1176
rect 4087 1162 4098 1170
rect 4148 1164 4155 1176
rect 4213 1170 4220 1176
rect 3927 1099 3929 1113
rect 3900 1076 3903 1082
rect 3877 1070 3903 1076
rect 3497 1064 3509 1070
rect 3537 1064 3549 1070
rect 3577 1064 3589 1070
rect 3617 1064 3629 1070
rect 3697 1064 3709 1070
rect 3737 1064 3749 1070
rect 3777 1064 3789 1070
rect 3817 1064 3829 1070
rect 3197 978 3209 984
rect 3237 978 3249 984
rect 3277 978 3289 984
rect 3349 978 3361 984
rect 3419 978 3431 984
rect 3477 978 3489 984
rect 3517 978 3529 984
rect 3557 978 3569 984
rect 3597 978 3609 984
rect 3637 978 3649 984
rect 3877 1024 3885 1070
rect 3921 1064 3929 1099
rect 3977 1093 3985 1142
rect 4037 1141 4045 1156
rect 4148 1157 4169 1164
rect 4127 1146 4133 1148
rect 4194 1146 4201 1152
rect 4037 1127 4053 1141
rect 4127 1140 4201 1146
rect 3977 1024 3985 1079
rect 4037 1064 4045 1127
rect 4053 1113 4067 1127
rect 4059 1068 4073 1076
rect 4127 1068 4133 1140
rect 4194 1132 4201 1140
rect 4206 1124 4240 1132
rect 4234 1119 4240 1124
rect 4187 1106 4214 1113
rect 4093 1062 4133 1068
rect 4141 1068 4185 1074
rect 4093 1044 4099 1062
rect 4141 1054 4147 1068
rect 4253 1072 4259 1156
rect 4309 1148 4321 1156
rect 4369 1156 4397 1162
rect 4357 1153 4409 1156
rect 4549 1156 4577 1162
rect 4297 1142 4321 1148
rect 4417 1142 4425 1156
rect 4479 1148 4491 1156
rect 4537 1153 4589 1156
rect 4479 1142 4503 1148
rect 4597 1142 4605 1156
rect 4297 1093 4305 1142
rect 4400 1135 4425 1142
rect 4399 1113 4407 1135
rect 4197 1064 4259 1072
rect 4117 1048 4147 1054
rect 4165 1050 4203 1058
rect 4195 1044 4203 1050
rect 4087 1004 4099 1038
rect 4145 1030 4167 1042
rect 4195 1030 4213 1044
rect 4141 1024 4153 1030
rect 4195 1024 4203 1030
rect 4297 1024 4305 1079
rect 4393 1064 4401 1099
rect 4495 1093 4503 1142
rect 4580 1135 4605 1142
rect 4686 1138 4704 1140
rect 4579 1113 4587 1135
rect 4674 1129 4704 1138
rect 4696 1101 4704 1129
rect 3677 978 3689 984
rect 3717 978 3729 984
rect 3757 978 3769 984
rect 3797 978 3809 984
rect 3837 978 3849 984
rect 3899 978 3911 984
rect 3957 978 3969 984
rect 3997 978 4009 984
rect 4057 978 4069 984
rect 4115 978 4127 984
rect 4161 978 4173 984
rect 4227 978 4239 984
rect 4277 978 4289 984
rect 4317 978 4329 984
rect 4495 1024 4503 1079
rect 4573 1064 4581 1099
rect 4362 978 4374 984
rect 4412 978 4424 984
rect 4471 978 4483 984
rect 4511 978 4523 984
rect 4698 1032 4705 1087
rect 4658 1026 4705 1032
rect 4658 1024 4669 1026
rect 4542 978 4554 984
rect 4592 978 4604 984
rect 4697 1024 4705 1026
rect 4637 978 4649 984
rect 4677 978 4689 984
rect -62 976 4776 978
rect -62 964 4 976
rect -62 962 4776 964
rect -62 498 -2 962
rect 31 956 43 962
rect 71 956 83 962
rect 127 956 139 962
rect 171 956 183 962
rect 55 861 63 916
rect 216 956 228 962
rect 266 956 278 962
rect 371 956 383 962
rect 449 956 461 962
rect 497 956 509 962
rect 591 956 603 962
rect 671 956 683 962
rect 717 956 729 962
rect 757 956 769 962
rect 847 956 859 962
rect 891 956 903 962
rect 55 798 63 847
rect 111 841 119 876
rect 111 827 113 841
rect 39 792 63 798
rect 39 784 51 792
rect 111 784 119 827
rect 154 802 162 916
rect 323 950 351 956
rect 363 878 391 884
rect 239 841 247 876
rect 332 870 344 876
rect 332 864 359 870
rect 353 841 359 864
rect 431 841 439 876
rect 475 870 483 916
rect 457 864 483 870
rect 457 858 460 864
rect 233 805 241 827
rect 145 794 183 802
rect 171 784 183 794
rect 215 798 240 805
rect 215 784 223 798
rect 111 774 121 784
rect 231 784 283 787
rect 360 784 367 827
rect 431 827 433 841
rect 431 784 439 827
rect 453 802 460 858
rect 516 833 524 916
rect 576 833 584 916
rect 738 914 749 916
rect 777 914 785 916
rect 738 908 785 914
rect 691 882 703 884
rect 663 876 703 882
rect 634 841 642 876
rect 778 853 785 908
rect 917 956 929 962
rect 957 956 969 962
rect 1031 956 1043 962
rect 1071 956 1083 962
rect 831 841 839 876
rect 457 796 460 802
rect 457 790 479 796
rect 243 778 271 784
rect 471 764 479 790
rect 516 764 524 819
rect 576 764 584 819
rect 634 784 642 827
rect 776 811 784 839
rect 634 773 660 784
rect 69 738 81 744
rect 141 738 153 744
rect 251 738 263 744
rect 332 738 344 744
rect 388 738 400 744
rect 449 738 461 744
rect 497 738 509 744
rect 591 738 603 744
rect 638 738 650 744
rect 688 738 700 744
rect 754 802 784 811
rect 766 800 784 802
rect 831 827 833 841
rect 831 784 839 827
rect 874 802 882 916
rect 937 861 945 916
rect 1015 914 1023 916
rect 1102 956 1114 962
rect 1152 956 1164 962
rect 1231 956 1243 962
rect 1271 956 1283 962
rect 1051 914 1062 916
rect 1015 908 1062 914
rect 1015 853 1022 908
rect 1215 914 1223 916
rect 1297 956 1309 962
rect 1362 956 1374 962
rect 1412 956 1424 962
rect 1251 914 1262 916
rect 1215 908 1262 914
rect 865 794 903 802
rect 891 784 903 794
rect 937 798 945 847
rect 1133 841 1141 876
rect 1215 853 1222 908
rect 1016 811 1024 839
rect 1016 802 1046 811
rect 1139 805 1147 827
rect 1216 811 1224 839
rect 1316 833 1324 916
rect 1471 956 1483 962
rect 1511 956 1523 962
rect 1537 956 1549 962
rect 1577 956 1589 962
rect 1636 956 1648 962
rect 1686 956 1698 962
rect 1393 841 1401 876
rect 1495 861 1503 916
rect 1557 861 1565 916
rect 1587 877 1603 883
rect 1597 867 1603 877
rect 1016 800 1034 802
rect 937 792 961 798
rect 949 784 961 792
rect 831 774 841 784
rect 1140 798 1165 805
rect 1216 802 1246 811
rect 1216 800 1234 802
rect 1097 784 1149 787
rect 1109 778 1137 784
rect 1157 784 1165 798
rect 1316 764 1324 819
rect 1399 805 1407 827
rect 1400 798 1425 805
rect 1495 798 1503 847
rect 1357 784 1409 787
rect 718 738 730 744
rect 861 738 873 744
rect 919 738 931 744
rect 1070 738 1082 744
rect 1117 738 1129 744
rect 1270 738 1282 744
rect 1369 778 1397 784
rect 1417 784 1425 798
rect 1479 792 1503 798
rect 1557 798 1565 847
rect 1617 823 1623 933
rect 1717 956 1729 962
rect 1761 956 1773 962
rect 1851 956 1863 962
rect 1659 841 1667 876
rect 1617 817 1633 823
rect 1653 805 1661 827
rect 1635 798 1660 805
rect 1738 802 1746 916
rect 1891 956 1903 962
rect 1931 956 1943 962
rect 1957 956 1969 962
rect 2051 956 2063 962
rect 2091 956 2103 962
rect 1781 841 1789 876
rect 1787 827 1789 841
rect 1836 833 1844 916
rect 1915 861 1923 916
rect 1557 792 1581 798
rect 1479 784 1491 792
rect 1569 784 1581 792
rect 1635 784 1643 798
rect 1717 794 1755 802
rect 1297 738 1309 744
rect 1377 738 1389 744
rect 1509 738 1521 744
rect 1651 784 1703 787
rect 1663 778 1691 784
rect 1717 784 1729 794
rect 1781 784 1789 827
rect 1779 774 1789 784
rect 1836 764 1844 819
rect 1915 798 1923 847
rect 1976 833 1984 916
rect 2035 914 2043 916
rect 2117 956 2129 962
rect 2182 956 2194 962
rect 2232 956 2244 962
rect 2331 956 2343 962
rect 2377 956 2389 962
rect 2437 956 2449 962
rect 2477 956 2489 962
rect 2571 956 2583 962
rect 2611 956 2623 962
rect 2657 956 2669 962
rect 2751 956 2763 962
rect 2791 956 2803 962
rect 2071 914 2082 916
rect 2035 908 2082 914
rect 2035 853 2042 908
rect 1899 792 1923 798
rect 1899 784 1911 792
rect 1976 764 1984 819
rect 2036 811 2044 839
rect 2136 833 2144 916
rect 2351 882 2363 884
rect 2323 876 2363 882
rect 2213 841 2221 876
rect 2294 841 2302 876
rect 2036 802 2066 811
rect 2396 833 2404 916
rect 2458 914 2469 916
rect 2497 914 2505 916
rect 2458 908 2505 914
rect 2498 853 2505 908
rect 2555 914 2563 916
rect 2591 914 2602 916
rect 2555 908 2602 914
rect 2555 853 2562 908
rect 2637 882 2649 884
rect 2637 876 2677 882
rect 2841 956 2853 962
rect 2911 956 2923 962
rect 2971 956 2983 962
rect 3051 956 3063 962
rect 3131 956 3143 962
rect 2698 841 2706 876
rect 2775 861 2783 916
rect 2036 800 2054 802
rect 1539 738 1551 744
rect 1671 738 1683 744
rect 1747 738 1759 744
rect 1851 738 1863 744
rect 1929 738 1941 744
rect 2136 764 2144 819
rect 2219 805 2227 827
rect 2220 798 2245 805
rect 2177 784 2229 787
rect 1957 738 1969 744
rect 2090 738 2102 744
rect 2189 778 2217 784
rect 2237 784 2245 798
rect 2294 784 2302 827
rect 2294 773 2320 784
rect 2396 764 2404 819
rect 2496 811 2504 839
rect 2117 738 2129 744
rect 2197 738 2209 744
rect 2298 738 2310 744
rect 2348 738 2360 744
rect 2474 802 2504 811
rect 2486 800 2504 802
rect 2556 811 2564 839
rect 2556 802 2586 811
rect 2556 800 2574 802
rect 2698 784 2706 827
rect 2775 798 2783 847
rect 2875 841 2883 876
rect 2876 801 2884 827
rect 2956 833 2964 916
rect 3157 956 3169 962
rect 3222 956 3234 962
rect 3272 956 3284 962
rect 3023 869 3040 876
rect 3103 869 3120 876
rect 3033 821 3040 869
rect 3113 821 3120 869
rect 3176 833 3184 916
rect 3317 956 3329 962
rect 3357 956 3369 962
rect 3417 956 3429 962
rect 3475 956 3487 962
rect 3521 956 3533 962
rect 3587 956 3599 962
rect 3659 956 3671 962
rect 3741 956 3753 962
rect 3807 956 3819 962
rect 3853 956 3865 962
rect 3911 956 3923 962
rect 3976 956 3988 962
rect 4026 956 4038 962
rect 4077 956 4089 962
rect 4135 956 4147 962
rect 4181 956 4193 962
rect 4247 956 4259 962
rect 4321 956 4333 962
rect 4387 956 4399 962
rect 4433 956 4445 962
rect 4491 956 4503 962
rect 4542 956 4554 962
rect 4592 956 4604 962
rect 3253 841 3261 876
rect 3337 861 3345 916
rect 3447 902 3459 936
rect 3501 910 3513 916
rect 3555 910 3563 916
rect 3505 898 3527 910
rect 3555 896 3573 910
rect 3453 878 3459 896
rect 3477 886 3507 892
rect 3555 890 3563 896
rect 2377 738 2389 744
rect 2438 738 2450 744
rect 2610 738 2622 744
rect 2680 773 2706 784
rect 2759 792 2783 798
rect 2855 794 2884 801
rect 2759 784 2771 792
rect 2855 784 2861 794
rect 2871 784 2923 786
rect 2843 744 2871 750
rect 2883 780 2911 784
rect 2956 764 2964 819
rect 3033 764 3040 807
rect 3113 764 3120 807
rect 3176 764 3184 819
rect 3259 805 3267 827
rect 3260 798 3285 805
rect 3217 784 3269 787
rect 2640 738 2652 744
rect 2690 738 2702 744
rect 2789 738 2801 744
rect 2891 738 2903 744
rect 2971 738 2983 744
rect 3011 738 3023 744
rect 3051 738 3063 744
rect 3091 738 3103 744
rect 3131 738 3143 744
rect 3229 778 3257 784
rect 3277 784 3285 798
rect 3337 798 3345 847
rect 3397 813 3405 876
rect 3419 864 3433 872
rect 3453 872 3493 878
rect 3413 813 3427 827
rect 3397 799 3413 813
rect 3487 800 3493 872
rect 3501 872 3507 886
rect 3525 882 3563 890
rect 3501 866 3545 872
rect 3557 868 3619 876
rect 3547 827 3574 834
rect 3594 816 3600 821
rect 3566 808 3600 816
rect 3554 800 3561 808
rect 3337 792 3361 798
rect 3349 784 3361 792
rect 3397 784 3405 799
rect 3487 794 3561 800
rect 3487 792 3493 794
rect 3554 788 3561 794
rect 3447 770 3458 778
rect 3451 764 3458 770
rect 3508 776 3529 783
rect 3613 784 3619 868
rect 3637 870 3645 916
rect 3777 910 3785 916
rect 3827 910 3839 916
rect 3767 896 3785 910
rect 3813 898 3835 910
rect 3881 902 3893 936
rect 3777 890 3785 896
rect 3777 882 3815 890
rect 3833 886 3863 892
rect 3637 864 3663 870
rect 3660 858 3663 864
rect 3660 802 3667 858
rect 3681 841 3689 876
rect 3687 827 3689 841
rect 3660 796 3663 802
rect 3508 764 3515 776
rect 3573 764 3580 770
rect 3567 758 3580 764
rect 3641 790 3663 796
rect 3641 764 3649 790
rect 3681 784 3689 827
rect 3721 868 3783 876
rect 3721 784 3727 868
rect 3833 872 3839 886
rect 3881 878 3887 896
rect 3795 866 3839 872
rect 3847 872 3887 878
rect 3766 827 3793 834
rect 3740 816 3746 821
rect 3740 808 3774 816
rect 3779 800 3786 808
rect 3847 800 3853 872
rect 4107 902 4119 936
rect 4161 910 4173 916
rect 4215 910 4223 916
rect 4165 898 4187 910
rect 4215 896 4233 910
rect 4113 878 4119 896
rect 4137 886 4167 892
rect 4215 890 4223 896
rect 3907 864 3921 872
rect 3913 813 3927 827
rect 3935 813 3943 876
rect 3999 841 4007 876
rect 3779 794 3853 800
rect 3927 799 3943 813
rect 3993 805 4001 827
rect 4057 813 4065 876
rect 4079 864 4093 872
rect 4113 872 4153 878
rect 4073 813 4087 827
rect 3779 788 3786 794
rect 3847 792 3853 794
rect 3811 776 3832 783
rect 3935 784 3943 799
rect 3975 798 4000 805
rect 4057 799 4073 813
rect 4147 800 4153 872
rect 4161 872 4167 886
rect 4185 882 4223 890
rect 4161 866 4205 872
rect 4217 868 4279 876
rect 4207 827 4234 834
rect 4254 816 4260 821
rect 4226 808 4260 816
rect 4214 800 4221 808
rect 3975 784 3983 798
rect 3760 764 3767 770
rect 3825 764 3832 776
rect 3882 770 3893 778
rect 3882 764 3889 770
rect 3760 758 3773 764
rect 3991 784 4043 787
rect 4003 778 4031 784
rect 4057 784 4065 799
rect 4147 794 4221 800
rect 4147 792 4153 794
rect 4214 788 4221 794
rect 4107 770 4118 778
rect 4111 764 4118 770
rect 4168 776 4189 783
rect 4273 784 4279 868
rect 4168 764 4175 776
rect 4233 764 4240 770
rect 4227 758 4240 764
rect 4357 910 4365 916
rect 4407 910 4419 916
rect 4347 896 4365 910
rect 4393 898 4415 910
rect 4461 902 4473 936
rect 4357 890 4365 896
rect 4357 882 4395 890
rect 4413 886 4443 892
rect 4301 868 4363 876
rect 4301 784 4307 868
rect 4413 872 4419 886
rect 4461 878 4467 896
rect 4375 866 4419 872
rect 4427 872 4467 878
rect 4346 827 4373 834
rect 4320 816 4326 821
rect 4320 808 4354 816
rect 4359 800 4366 808
rect 4427 800 4433 872
rect 4642 956 4654 962
rect 4692 956 4704 962
rect 4487 864 4501 872
rect 4493 813 4507 827
rect 4515 813 4523 876
rect 4573 841 4581 876
rect 4673 841 4681 876
rect 4359 794 4433 800
rect 4507 799 4523 813
rect 4579 805 4587 827
rect 4679 805 4687 827
rect 4359 788 4366 794
rect 4427 792 4433 794
rect 4391 776 4412 783
rect 4515 784 4523 799
rect 4580 798 4605 805
rect 4680 798 4705 805
rect 4340 764 4347 770
rect 4405 764 4412 776
rect 4462 770 4473 778
rect 4462 764 4469 770
rect 4340 758 4353 764
rect 4537 784 4589 787
rect 4549 778 4577 784
rect 4597 784 4605 798
rect 4637 784 4689 787
rect 4649 778 4677 784
rect 4697 784 4705 798
rect 3157 738 3169 744
rect 3237 738 3249 744
rect 3319 738 3331 744
rect 3419 738 3431 744
rect 3477 738 3489 744
rect 3525 738 3537 744
rect 3587 738 3599 744
rect 3659 738 3671 744
rect 3741 738 3753 744
rect 3803 738 3815 744
rect 3851 738 3863 744
rect 3909 738 3921 744
rect 4011 738 4023 744
rect 4079 738 4091 744
rect 4137 738 4149 744
rect 4185 738 4197 744
rect 4247 738 4259 744
rect 4321 738 4333 744
rect 4383 738 4395 744
rect 4431 738 4443 744
rect 4489 738 4501 744
rect 4557 738 4569 744
rect 4657 738 4669 744
rect 4782 738 4842 1202
rect 4 736 4842 738
rect 4776 724 4842 736
rect 4 722 4842 724
rect 31 716 43 722
rect 71 716 83 722
rect 118 716 130 722
rect 168 716 180 722
rect 53 653 60 696
rect 114 676 140 687
rect 197 716 209 722
rect 278 716 290 722
rect 328 716 340 722
rect 53 591 60 639
rect 114 633 122 676
rect 216 641 224 696
rect 274 676 300 687
rect 358 716 370 722
rect 511 716 523 722
rect 589 716 601 722
rect 691 716 703 722
rect 769 716 781 722
rect 847 716 859 722
rect 937 716 949 722
rect 1071 716 1083 722
rect 1151 716 1163 722
rect 274 633 282 676
rect 475 662 483 676
rect 503 676 531 682
rect 491 673 543 676
rect 406 658 424 660
rect 43 584 60 591
rect 114 584 122 619
rect 143 578 183 584
rect 171 576 183 578
rect 216 544 224 627
rect 394 649 424 658
rect 475 655 500 662
rect 416 621 424 649
rect 493 633 501 655
rect 274 584 282 619
rect 571 633 579 676
rect 611 670 619 696
rect 597 664 619 670
rect 597 658 600 664
rect 571 619 573 633
rect 303 578 343 584
rect 331 576 343 578
rect 418 552 425 607
rect 499 584 507 619
rect 571 584 579 619
rect 593 602 600 658
rect 655 662 663 676
rect 683 676 711 682
rect 671 673 723 676
rect 655 655 680 662
rect 673 633 681 655
rect 751 633 759 676
rect 791 670 799 696
rect 777 664 799 670
rect 879 676 889 686
rect 817 666 829 676
rect 777 658 780 664
rect 817 658 855 666
rect 751 619 753 633
rect 597 596 600 602
rect 597 590 623 596
rect 378 546 425 552
rect 378 544 389 546
rect 417 544 425 546
rect 615 544 623 590
rect 679 584 687 619
rect 751 584 759 619
rect 773 602 780 658
rect 777 596 780 602
rect 777 590 803 596
rect 795 544 803 590
rect 838 544 846 658
rect 881 633 889 676
rect 929 676 957 682
rect 917 673 969 676
rect 977 662 985 676
rect 960 655 985 662
rect 1035 662 1043 676
rect 1063 676 1091 682
rect 1180 716 1192 722
rect 1230 716 1242 722
rect 1311 716 1323 722
rect 1357 716 1369 722
rect 1457 716 1469 722
rect 1558 716 1570 722
rect 1608 716 1620 722
rect 1220 676 1246 687
rect 1051 673 1103 676
rect 1035 655 1060 662
rect 887 619 889 633
rect 959 633 967 655
rect 1053 633 1061 655
rect 1136 633 1144 676
rect 1238 633 1246 676
rect 1296 641 1304 696
rect 1349 676 1377 682
rect 1337 673 1389 676
rect 1449 676 1477 682
rect 1397 662 1405 676
rect 1437 673 1489 676
rect 1554 676 1580 687
rect 1640 716 1652 722
rect 1690 716 1702 722
rect 1738 716 1750 722
rect 1857 716 1869 722
rect 1958 716 1970 722
rect 2008 716 2020 722
rect 2057 716 2069 722
rect 2210 716 2222 722
rect 2291 716 2303 722
rect 2357 716 2369 722
rect 2438 716 2450 722
rect 2538 716 2550 722
rect 2671 716 2683 722
rect 1680 676 1706 687
rect 1497 662 1505 676
rect 1380 655 1405 662
rect 1480 655 1505 662
rect 881 584 889 619
rect 953 584 961 619
rect 1059 584 1067 619
rect 1136 584 1144 619
rect 1238 584 1246 619
rect 71 498 83 504
rect 151 498 163 504
rect 197 498 209 504
rect 311 498 323 504
rect 357 498 369 504
rect 397 498 409 504
rect 476 498 488 504
rect 526 498 538 504
rect 589 498 601 504
rect 656 498 668 504
rect 706 498 718 504
rect 769 498 781 504
rect 817 498 829 504
rect 861 498 873 504
rect 922 498 934 504
rect 972 498 984 504
rect 1177 578 1217 584
rect 1177 576 1189 578
rect 1296 544 1304 627
rect 1379 633 1387 655
rect 1479 633 1487 655
rect 1554 633 1562 676
rect 1698 633 1706 676
rect 1849 676 1877 682
rect 1837 673 1889 676
rect 1954 676 1980 687
rect 2049 676 2077 682
rect 1897 662 1905 676
rect 1786 658 1804 660
rect 1774 649 1804 658
rect 1880 655 1905 662
rect 1796 621 1804 649
rect 1373 584 1381 619
rect 1473 584 1481 619
rect 1554 584 1562 619
rect 1698 584 1706 619
rect 1879 633 1887 655
rect 1907 637 1923 643
rect 1036 498 1048 504
rect 1086 498 1098 504
rect 1151 498 1163 504
rect 1197 498 1209 504
rect 1311 498 1323 504
rect 1342 498 1354 504
rect 1392 498 1404 504
rect 1583 578 1623 584
rect 1611 576 1623 578
rect 1637 578 1677 584
rect 1637 576 1649 578
rect 1798 552 1805 607
rect 1873 584 1881 619
rect 1758 546 1805 552
rect 1758 544 1769 546
rect 1797 544 1805 546
rect 1917 563 1923 637
rect 1954 633 1962 676
rect 2037 673 2089 676
rect 2137 677 2153 683
rect 2097 662 2105 676
rect 2137 663 2143 677
rect 2080 655 2105 662
rect 2117 657 2143 663
rect 2156 658 2174 660
rect 2079 633 2087 655
rect 1954 584 1962 619
rect 2073 584 2081 619
rect 2117 587 2123 657
rect 2156 649 2186 658
rect 2255 662 2263 676
rect 2283 676 2311 682
rect 2271 673 2323 676
rect 2349 676 2377 682
rect 2337 673 2389 676
rect 2397 662 2405 676
rect 2255 655 2280 662
rect 2380 655 2405 662
rect 2486 658 2504 660
rect 2156 621 2164 649
rect 2273 633 2281 655
rect 1907 557 1923 563
rect 1983 578 2023 584
rect 2011 576 2023 578
rect 2155 552 2162 607
rect 2237 563 2243 633
rect 2379 633 2387 655
rect 2474 649 2504 658
rect 2698 716 2710 722
rect 2821 716 2833 722
rect 2883 716 2895 722
rect 2931 716 2943 722
rect 2989 716 3001 722
rect 3057 716 3069 722
rect 3137 716 3149 722
rect 3197 716 3209 722
rect 3258 716 3270 722
rect 3391 716 3403 722
rect 3469 716 3481 722
rect 3551 716 3563 722
rect 3621 716 3633 722
rect 3683 716 3695 722
rect 3731 716 3743 722
rect 3789 716 3801 722
rect 3857 716 3869 722
rect 3989 716 4001 722
rect 4039 716 4051 722
rect 4097 716 4109 722
rect 4145 716 4157 722
rect 4207 716 4219 722
rect 4259 716 4271 722
rect 4339 716 4351 722
rect 4471 716 4483 722
rect 4541 716 4553 722
rect 4603 716 4615 722
rect 4651 716 4663 722
rect 4709 716 4721 722
rect 2586 658 2604 660
rect 2574 649 2604 658
rect 2496 621 2504 649
rect 2596 621 2604 649
rect 2656 641 2664 696
rect 2840 696 2853 702
rect 2840 690 2847 696
rect 2905 684 2912 696
rect 2746 658 2764 660
rect 2734 649 2764 658
rect 2279 584 2287 619
rect 2373 584 2381 619
rect 2227 557 2243 563
rect 2155 546 2202 552
rect 2155 544 2163 546
rect 2191 544 2202 546
rect 1442 498 1454 504
rect 1492 498 1504 504
rect 1591 498 1603 504
rect 1657 498 1669 504
rect 1737 498 1749 504
rect 1777 498 1789 504
rect 1842 498 1854 504
rect 1892 498 1904 504
rect 1991 498 2003 504
rect 2042 498 2054 504
rect 2092 498 2104 504
rect 2171 498 2183 504
rect 2211 498 2223 504
rect 2256 498 2268 504
rect 2306 498 2318 504
rect 2498 552 2505 607
rect 2598 552 2605 607
rect 2458 546 2505 552
rect 2458 544 2469 546
rect 2342 498 2354 504
rect 2392 498 2404 504
rect 2497 544 2505 546
rect 2558 546 2605 552
rect 2558 544 2569 546
rect 2597 544 2605 546
rect 2656 544 2664 627
rect 2756 621 2764 649
rect 2758 552 2765 607
rect 2718 546 2765 552
rect 2718 544 2729 546
rect 2437 498 2449 504
rect 2477 498 2489 504
rect 2537 498 2549 504
rect 2577 498 2589 504
rect 2671 498 2683 504
rect 2757 544 2765 546
rect 2801 592 2807 676
rect 2891 677 2912 684
rect 2962 690 2969 696
rect 2962 682 2973 690
rect 2859 666 2866 672
rect 2927 666 2933 668
rect 2859 660 2933 666
rect 3015 661 3023 676
rect 3049 676 3077 682
rect 3037 673 3089 676
rect 3097 662 3105 676
rect 2859 652 2866 660
rect 2820 644 2854 652
rect 2820 639 2826 644
rect 2846 626 2873 633
rect 2801 584 2863 592
rect 2875 588 2919 594
rect 2857 570 2895 578
rect 2913 574 2919 588
rect 2927 588 2933 660
rect 3007 647 3023 661
rect 3080 655 3105 662
rect 2993 633 3007 647
rect 2927 582 2967 588
rect 2987 588 3001 596
rect 3015 584 3023 647
rect 3079 633 3087 655
rect 3156 641 3164 696
rect 3216 641 3224 696
rect 3306 658 3324 660
rect 3294 649 3324 658
rect 3073 584 3081 619
rect 2857 564 2865 570
rect 2913 568 2943 574
rect 2961 564 2967 582
rect 2847 550 2865 564
rect 2893 550 2915 562
rect 2857 544 2865 550
rect 2907 544 2919 550
rect 2961 524 2973 558
rect 3156 544 3164 627
rect 3216 544 3224 627
rect 3316 621 3324 649
rect 3376 641 3384 696
rect 3439 668 3451 676
rect 3439 662 3463 668
rect 3318 552 3325 607
rect 3278 546 3325 552
rect 3278 544 3289 546
rect 2697 498 2709 504
rect 2737 498 2749 504
rect 2821 498 2833 504
rect 2887 498 2899 504
rect 2933 498 2945 504
rect 2991 498 3003 504
rect 3042 498 3054 504
rect 3092 498 3104 504
rect 3317 544 3325 546
rect 3376 544 3384 627
rect 3455 613 3463 662
rect 3515 662 3523 676
rect 3543 676 3571 682
rect 3531 673 3583 676
rect 3640 696 3653 702
rect 3640 690 3647 696
rect 3705 684 3712 696
rect 3515 655 3540 662
rect 3533 633 3541 655
rect 3455 544 3463 599
rect 3539 584 3547 619
rect 3601 592 3607 676
rect 3691 677 3712 684
rect 3762 690 3769 696
rect 3762 682 3773 690
rect 3659 666 3666 672
rect 3727 666 3733 668
rect 3659 660 3733 666
rect 3815 661 3823 676
rect 3849 676 3877 682
rect 3837 673 3889 676
rect 4187 696 4200 702
rect 4071 690 4078 696
rect 4067 682 4078 690
rect 4128 684 4135 696
rect 4193 690 4200 696
rect 3897 662 3905 676
rect 3959 668 3971 676
rect 3959 662 3983 668
rect 3659 652 3666 660
rect 3620 644 3654 652
rect 3620 639 3626 644
rect 3646 626 3673 633
rect 3601 584 3663 592
rect 3675 588 3719 594
rect 3137 498 3149 504
rect 3197 498 3209 504
rect 3257 498 3269 504
rect 3297 498 3309 504
rect 3391 498 3403 504
rect 3431 498 3443 504
rect 3471 498 3483 504
rect 3657 570 3695 578
rect 3713 574 3719 588
rect 3727 588 3733 660
rect 3807 647 3823 661
rect 3880 655 3905 662
rect 3793 633 3807 647
rect 3727 582 3767 588
rect 3787 588 3801 596
rect 3815 584 3823 647
rect 3879 633 3887 655
rect 3873 584 3881 619
rect 3975 613 3983 662
rect 4017 661 4025 676
rect 4128 677 4149 684
rect 4107 666 4113 668
rect 4174 666 4181 672
rect 4017 647 4033 661
rect 4107 660 4181 666
rect 3657 564 3665 570
rect 3713 568 3743 574
rect 3761 564 3767 582
rect 3647 550 3665 564
rect 3693 550 3715 562
rect 3657 544 3665 550
rect 3707 544 3719 550
rect 3761 524 3773 558
rect 3975 544 3983 599
rect 4017 584 4025 647
rect 4033 633 4047 647
rect 4039 588 4053 596
rect 3516 498 3528 504
rect 3566 498 3578 504
rect 3621 498 3633 504
rect 3687 498 3699 504
rect 3733 498 3745 504
rect 3791 498 3803 504
rect 3842 498 3854 504
rect 3892 498 3904 504
rect 4107 588 4113 660
rect 4174 652 4181 660
rect 4186 644 4220 652
rect 4214 639 4220 644
rect 4167 626 4194 633
rect 4073 582 4113 588
rect 4121 588 4165 594
rect 4073 564 4079 582
rect 4121 574 4127 588
rect 4233 592 4239 676
rect 4289 668 4301 676
rect 4369 668 4381 676
rect 4277 662 4301 668
rect 4357 662 4381 668
rect 4435 662 4443 676
rect 4463 676 4491 682
rect 4451 673 4503 676
rect 4560 696 4573 702
rect 4560 690 4567 696
rect 4625 684 4632 696
rect 4277 613 4285 662
rect 4357 613 4365 662
rect 4435 655 4460 662
rect 4453 633 4461 655
rect 4177 584 4239 592
rect 4097 568 4127 574
rect 4145 570 4183 578
rect 4175 564 4183 570
rect 4067 524 4079 558
rect 4125 550 4147 562
rect 4175 550 4193 564
rect 4121 544 4133 550
rect 4175 544 4183 550
rect 4277 544 4285 599
rect 4357 544 4365 599
rect 4459 584 4467 619
rect 4521 592 4527 676
rect 4611 677 4632 684
rect 4682 690 4689 696
rect 4682 682 4693 690
rect 4579 666 4586 672
rect 4647 666 4653 668
rect 4579 660 4653 666
rect 4735 661 4743 676
rect 4579 652 4586 660
rect 4540 644 4574 652
rect 4540 639 4546 644
rect 4566 626 4593 633
rect 4521 584 4583 592
rect 4595 588 4639 594
rect 3951 498 3963 504
rect 3991 498 4003 504
rect 4037 498 4049 504
rect 4095 498 4107 504
rect 4141 498 4153 504
rect 4207 498 4219 504
rect 4257 498 4269 504
rect 4297 498 4309 504
rect 4337 498 4349 504
rect 4377 498 4389 504
rect 4577 570 4615 578
rect 4633 574 4639 588
rect 4647 588 4653 660
rect 4727 647 4743 661
rect 4713 633 4727 647
rect 4647 582 4687 588
rect 4707 588 4721 596
rect 4735 584 4743 647
rect 4577 564 4585 570
rect 4633 568 4663 574
rect 4681 564 4687 582
rect 4567 550 4585 564
rect 4613 550 4635 562
rect 4577 544 4585 550
rect 4627 544 4639 550
rect 4681 524 4693 558
rect 4436 498 4448 504
rect 4486 498 4498 504
rect 4541 498 4553 504
rect 4607 498 4619 504
rect 4653 498 4665 504
rect 4711 498 4723 504
rect -62 496 4776 498
rect -62 484 4 496
rect -62 482 4776 484
rect -62 18 -2 482
rect 17 476 29 482
rect 57 476 69 482
rect 97 476 109 482
rect 137 476 149 482
rect 191 476 203 482
rect 231 476 243 482
rect 271 476 283 482
rect 311 476 323 482
rect 367 476 379 482
rect 411 476 423 482
rect 37 381 45 436
rect 117 381 125 436
rect 215 381 223 436
rect 247 397 263 403
rect 37 318 45 367
rect 117 318 125 367
rect 215 318 223 367
rect 257 347 263 397
rect 295 381 303 436
rect 451 476 463 482
rect 491 476 503 482
rect 551 476 563 482
rect 591 476 603 482
rect 691 476 703 482
rect 791 476 803 482
rect 295 318 303 367
rect 351 361 359 396
rect 351 347 353 361
rect 37 312 61 318
rect 117 312 141 318
rect 49 304 61 312
rect 129 304 141 312
rect 199 312 223 318
rect 279 312 303 318
rect 199 304 211 312
rect 279 304 291 312
rect 351 304 359 347
rect 394 322 402 436
rect 427 397 443 403
rect 385 314 423 322
rect 411 304 423 314
rect 437 307 443 397
rect 475 381 483 436
rect 535 434 543 436
rect 571 434 582 436
rect 535 428 582 434
rect 535 373 542 428
rect 643 470 671 476
rect 683 398 711 404
rect 831 476 843 482
rect 871 476 883 482
rect 897 476 909 482
rect 937 476 949 482
rect 991 476 1003 482
rect 1031 476 1043 482
rect 1071 476 1083 482
rect 1111 476 1123 482
rect 1211 476 1223 482
rect 1262 476 1274 482
rect 1312 476 1324 482
rect 1411 476 1423 482
rect 652 390 664 396
rect 652 384 679 390
rect 763 389 780 396
rect 475 318 483 367
rect 673 361 679 384
rect 536 331 544 359
rect 536 322 566 331
rect 536 320 554 322
rect 459 312 483 318
rect 351 294 361 304
rect 459 304 471 312
rect 680 304 687 347
rect 773 341 780 389
rect 855 381 863 436
rect 917 381 925 436
rect 1015 381 1023 436
rect 1095 381 1103 436
rect 1163 470 1191 476
rect 1203 398 1231 404
rect 1442 476 1454 482
rect 1492 476 1504 482
rect 1537 476 1549 482
rect 1651 476 1663 482
rect 1697 476 1709 482
rect 1757 476 1769 482
rect 1797 476 1809 482
rect 1877 476 1889 482
rect 1957 476 1969 482
rect 1997 476 2009 482
rect 1172 390 1184 396
rect 1172 384 1199 390
rect 19 258 31 264
rect 99 258 111 264
rect 229 258 241 264
rect 309 258 321 264
rect 381 258 393 264
rect 489 258 501 264
rect 590 258 602 264
rect 773 284 780 327
rect 855 318 863 367
rect 839 312 863 318
rect 917 318 925 367
rect 1015 318 1023 367
rect 1095 318 1103 367
rect 1193 361 1199 384
rect 1293 361 1301 396
rect 1383 389 1400 396
rect 917 312 941 318
rect 839 304 851 312
rect 929 304 941 312
rect 652 258 664 264
rect 708 258 720 264
rect 751 258 763 264
rect 791 258 803 264
rect 869 258 881 264
rect 999 312 1023 318
rect 1079 312 1103 318
rect 999 304 1011 312
rect 1079 304 1091 312
rect 1200 304 1207 347
rect 1299 325 1307 347
rect 1393 341 1400 389
rect 1473 361 1481 396
rect 1556 353 1564 436
rect 1671 402 1683 404
rect 1643 396 1683 402
rect 1614 361 1622 396
rect 1300 318 1325 325
rect 1257 304 1309 307
rect 899 258 911 264
rect 1029 258 1041 264
rect 1109 258 1121 264
rect 1269 298 1297 304
rect 1317 304 1325 318
rect 1393 284 1400 327
rect 1479 325 1487 347
rect 1716 353 1724 436
rect 1778 434 1789 436
rect 1817 434 1825 436
rect 1778 428 1825 434
rect 1818 373 1825 428
rect 1857 402 1869 404
rect 1857 396 1897 402
rect 2037 476 2049 482
rect 2077 476 2089 482
rect 2117 476 2129 482
rect 2157 476 2169 482
rect 2251 476 2263 482
rect 1918 361 1926 396
rect 1977 381 1985 436
rect 1480 318 1505 325
rect 1437 304 1489 307
rect 1449 298 1477 304
rect 1497 304 1505 318
rect 1556 284 1564 339
rect 1614 304 1622 347
rect 1737 343 1743 353
rect 1614 293 1640 304
rect 1716 284 1724 339
rect 1737 337 1753 343
rect 1816 331 1824 359
rect 1172 258 1184 264
rect 1228 258 1240 264
rect 1277 258 1289 264
rect 1371 258 1383 264
rect 1411 258 1423 264
rect 1457 258 1469 264
rect 1537 258 1549 264
rect 1618 258 1630 264
rect 1668 258 1680 264
rect 1794 322 1824 331
rect 2057 381 2065 436
rect 1806 320 1824 322
rect 1918 304 1926 347
rect 1977 318 1985 367
rect 2017 323 2023 373
rect 1977 312 2001 318
rect 2017 317 2033 323
rect 2057 318 2065 367
rect 2097 327 2103 393
rect 2137 381 2145 436
rect 2187 397 2203 403
rect 2057 312 2081 318
rect 2137 318 2145 367
rect 2197 347 2203 397
rect 2291 476 2303 482
rect 2331 476 2343 482
rect 2357 476 2369 482
rect 2437 476 2449 482
rect 2477 476 2489 482
rect 2571 476 2583 482
rect 2631 476 2643 482
rect 2671 476 2683 482
rect 2717 476 2729 482
rect 2797 476 2809 482
rect 2891 476 2903 482
rect 2931 476 2943 482
rect 2223 389 2240 396
rect 2233 341 2240 389
rect 2315 381 2323 436
rect 2458 434 2469 436
rect 2497 434 2505 436
rect 2458 428 2505 434
rect 2380 389 2397 396
rect 2137 312 2161 318
rect 1989 304 2001 312
rect 2069 304 2081 312
rect 2149 304 2161 312
rect 1900 293 1926 304
rect 1697 258 1709 264
rect 1758 258 1770 264
rect 1860 258 1872 264
rect 1910 258 1922 264
rect 2233 284 2240 327
rect 2315 318 2323 367
rect 2380 341 2387 389
rect 2498 373 2505 428
rect 2496 331 2504 359
rect 2556 353 2564 436
rect 2615 434 2623 436
rect 2651 434 2662 436
rect 2615 428 2662 434
rect 2615 373 2622 428
rect 2697 402 2709 404
rect 2697 396 2737 402
rect 2976 476 2988 482
rect 3026 476 3038 482
rect 2758 361 2766 396
rect 2820 389 2837 396
rect 2299 312 2323 318
rect 2299 304 2311 312
rect 2380 284 2387 327
rect 1959 258 1971 264
rect 2039 258 2051 264
rect 2119 258 2131 264
rect 2211 258 2223 264
rect 2251 258 2263 264
rect 2329 258 2341 264
rect 2357 258 2369 264
rect 2397 258 2409 264
rect 2474 322 2504 331
rect 2486 320 2504 322
rect 2556 284 2564 339
rect 2616 331 2624 359
rect 2616 322 2646 331
rect 2616 320 2634 322
rect 2758 304 2766 347
rect 2820 341 2827 389
rect 2915 381 2923 436
rect 3076 476 3088 482
rect 3126 476 3138 482
rect 3211 476 3223 482
rect 3271 476 3283 482
rect 3316 476 3328 482
rect 3366 476 3378 482
rect 3451 476 3463 482
rect 3551 476 3563 482
rect 3607 476 3619 482
rect 3677 476 3689 482
rect 3717 476 3729 482
rect 2438 258 2450 264
rect 2571 258 2583 264
rect 2670 258 2682 264
rect 2740 293 2766 304
rect 2820 284 2827 327
rect 2915 318 2923 367
rect 2999 361 3007 396
rect 3099 361 3107 396
rect 3183 389 3200 396
rect 2993 325 3001 347
rect 3093 325 3101 347
rect 3193 341 3200 389
rect 3256 353 3264 436
rect 3471 402 3483 404
rect 3443 396 3483 402
rect 3757 476 3769 482
rect 3797 476 3809 482
rect 3856 476 3868 482
rect 3906 476 3918 482
rect 3971 476 3983 482
rect 4031 476 4043 482
rect 4077 476 4089 482
rect 4135 476 4147 482
rect 4181 476 4193 482
rect 4247 476 4259 482
rect 4311 476 4323 482
rect 4351 476 4363 482
rect 3639 397 3643 406
rect 3339 361 3347 396
rect 3414 361 3422 396
rect 3523 389 3540 396
rect 2899 312 2923 318
rect 2975 318 3000 325
rect 3075 318 3100 325
rect 2899 304 2911 312
rect 2975 304 2983 318
rect 2700 258 2712 264
rect 2750 258 2762 264
rect 2991 304 3043 307
rect 3075 304 3083 318
rect 3003 298 3031 304
rect 3091 304 3143 307
rect 3103 298 3131 304
rect 3193 284 3200 327
rect 3256 284 3264 339
rect 3333 325 3341 347
rect 3315 318 3340 325
rect 3315 304 3323 318
rect 3331 304 3383 307
rect 3343 298 3371 304
rect 3414 304 3422 347
rect 3533 341 3540 389
rect 3577 388 3585 396
rect 3577 380 3613 388
rect 3414 293 3440 304
rect 3533 284 3540 327
rect 3618 324 3624 379
rect 3634 353 3643 397
rect 3697 381 3705 436
rect 3777 381 3785 436
rect 3603 312 3613 318
rect 3603 284 3609 312
rect 3640 304 3647 339
rect 3697 318 3705 367
rect 3777 318 3785 367
rect 3879 361 3887 396
rect 3873 325 3881 347
rect 3956 353 3964 436
rect 4016 353 4024 436
rect 4107 422 4119 456
rect 4161 430 4173 436
rect 4215 430 4223 436
rect 4165 418 4187 430
rect 4215 416 4233 430
rect 4113 398 4119 416
rect 4137 406 4167 412
rect 4215 410 4223 416
rect 3855 318 3880 325
rect 3697 312 3721 318
rect 3777 312 3801 318
rect 3709 304 3721 312
rect 3789 304 3801 312
rect 3855 304 3863 318
rect 2797 258 2809 264
rect 2837 258 2849 264
rect 2929 258 2941 264
rect 3011 258 3023 264
rect 3111 258 3123 264
rect 3171 258 3183 264
rect 3211 258 3223 264
rect 3271 258 3283 264
rect 3351 258 3363 264
rect 3418 258 3430 264
rect 3468 258 3480 264
rect 3511 258 3523 264
rect 3551 258 3563 264
rect 3871 304 3923 307
rect 3883 298 3911 304
rect 3956 284 3964 339
rect 4016 284 4024 339
rect 4057 333 4065 396
rect 4079 384 4093 392
rect 4113 392 4153 398
rect 4073 333 4087 347
rect 4057 319 4073 333
rect 4147 320 4153 392
rect 4161 392 4167 406
rect 4185 402 4223 410
rect 4396 476 4408 482
rect 4446 476 4458 482
rect 4511 476 4523 482
rect 4557 476 4569 482
rect 4615 476 4627 482
rect 4661 476 4673 482
rect 4727 476 4739 482
rect 4161 386 4205 392
rect 4217 388 4279 396
rect 4207 347 4234 354
rect 4254 336 4260 341
rect 4226 328 4260 336
rect 4214 320 4221 328
rect 4057 304 4065 319
rect 4147 314 4221 320
rect 4147 312 4153 314
rect 4214 308 4221 314
rect 4107 290 4118 298
rect 4111 284 4118 290
rect 4168 296 4189 303
rect 4273 304 4279 388
rect 4335 381 4343 436
rect 4335 318 4343 367
rect 4419 361 4427 396
rect 4413 325 4421 347
rect 4496 353 4504 436
rect 4587 422 4599 456
rect 4641 430 4653 436
rect 4695 430 4703 436
rect 4645 418 4667 430
rect 4695 416 4713 430
rect 4593 398 4599 416
rect 4617 406 4647 412
rect 4695 410 4703 416
rect 4168 284 4175 296
rect 4233 284 4240 290
rect 4227 278 4240 284
rect 4319 312 4343 318
rect 4395 318 4420 325
rect 4319 304 4331 312
rect 4395 304 4403 318
rect 4411 304 4463 307
rect 4423 298 4451 304
rect 4496 284 4504 339
rect 4537 333 4545 396
rect 4559 384 4573 392
rect 4593 392 4633 398
rect 4553 333 4567 347
rect 4537 319 4553 333
rect 4627 320 4633 392
rect 4641 392 4647 406
rect 4665 402 4703 410
rect 4641 386 4685 392
rect 4697 388 4759 396
rect 4687 347 4714 354
rect 4734 336 4740 341
rect 4706 328 4740 336
rect 4694 320 4701 328
rect 4537 304 4545 319
rect 4627 314 4701 320
rect 4627 312 4633 314
rect 4694 308 4701 314
rect 4587 290 4598 298
rect 4591 284 4598 290
rect 4648 296 4669 303
rect 4753 304 4759 388
rect 4648 284 4655 296
rect 4713 284 4720 290
rect 4707 278 4720 284
rect 3577 258 3585 264
rect 3617 258 3629 264
rect 3679 258 3691 264
rect 3759 258 3771 264
rect 3891 258 3903 264
rect 3971 258 3983 264
rect 4031 258 4043 264
rect 4079 258 4091 264
rect 4137 258 4149 264
rect 4185 258 4197 264
rect 4247 258 4259 264
rect 4349 258 4361 264
rect 4431 258 4443 264
rect 4511 258 4523 264
rect 4559 258 4571 264
rect 4617 258 4629 264
rect 4665 258 4677 264
rect 4727 258 4739 264
rect 4782 258 4842 722
rect 4 256 4842 258
rect 4776 244 4842 256
rect 4 242 4842 244
rect 90 236 102 242
rect 36 178 54 180
rect 36 169 66 178
rect 120 236 132 242
rect 170 236 182 242
rect 271 236 283 242
rect 337 236 349 242
rect 490 236 502 242
rect 160 196 186 207
rect 36 141 44 169
rect 178 153 186 196
rect 235 182 243 196
rect 263 196 291 202
rect 251 193 303 196
rect 329 196 357 202
rect 317 193 369 196
rect 377 182 385 196
rect 235 175 260 182
rect 360 175 385 182
rect 436 178 454 180
rect 253 153 261 175
rect 359 153 367 175
rect 436 169 466 178
rect 518 236 530 242
rect 620 236 632 242
rect 670 236 682 242
rect 738 236 750 242
rect 788 236 800 242
rect 660 196 686 207
rect 566 178 584 180
rect 554 169 584 178
rect 436 141 444 169
rect 576 141 584 169
rect 35 72 42 127
rect 178 104 186 139
rect 259 104 267 139
rect 353 104 361 139
rect 117 98 157 104
rect 117 96 129 98
rect 35 66 82 72
rect 35 64 43 66
rect 71 64 82 66
rect 51 18 63 24
rect 91 18 103 24
rect 137 18 149 24
rect 236 18 248 24
rect 286 18 298 24
rect 435 72 442 127
rect 578 72 585 127
rect 597 107 603 173
rect 678 153 686 196
rect 734 196 760 207
rect 817 236 829 242
rect 931 236 943 242
rect 1011 236 1023 242
rect 1057 236 1069 242
rect 1157 236 1169 242
rect 1238 236 1250 242
rect 1338 236 1350 242
rect 1458 236 1470 242
rect 1508 236 1520 242
rect 734 153 742 196
rect 836 161 844 216
rect 895 182 903 196
rect 923 196 951 202
rect 911 193 963 196
rect 895 175 920 182
rect 913 153 921 175
rect 678 104 686 139
rect 734 104 742 139
rect 617 98 657 104
rect 617 96 629 98
rect 435 66 482 72
rect 435 64 443 66
rect 471 64 482 66
rect 538 66 585 72
rect 538 64 549 66
rect 322 18 334 24
rect 372 18 384 24
rect 451 18 463 24
rect 491 18 503 24
rect 577 64 585 66
rect 763 98 803 104
rect 791 96 803 98
rect 836 64 844 147
rect 919 104 927 139
rect 977 127 983 193
rect 996 161 1004 216
rect 1049 196 1077 202
rect 1037 193 1089 196
rect 1149 196 1177 202
rect 1097 182 1105 196
rect 1137 193 1189 196
rect 1197 182 1205 196
rect 1080 175 1105 182
rect 1180 175 1205 182
rect 1286 178 1304 180
rect 996 64 1004 147
rect 1079 153 1087 175
rect 1179 153 1187 175
rect 1274 169 1304 178
rect 1454 196 1480 207
rect 1538 236 1550 242
rect 1658 236 1670 242
rect 1708 236 1720 242
rect 1386 178 1404 180
rect 1374 169 1404 178
rect 1296 141 1304 169
rect 1396 141 1404 169
rect 1454 153 1462 196
rect 1654 196 1680 207
rect 1738 236 1750 242
rect 1839 236 1851 242
rect 1939 236 1951 242
rect 2041 236 2053 242
rect 2119 236 2131 242
rect 2178 236 2190 242
rect 2280 236 2292 242
rect 2336 236 2348 242
rect 2417 236 2429 242
rect 2518 236 2530 242
rect 2568 236 2580 242
rect 2617 236 2629 242
rect 2697 236 2709 242
rect 2758 236 2770 242
rect 2857 236 2869 242
rect 2941 236 2953 242
rect 3003 236 3015 242
rect 3051 236 3063 242
rect 3109 236 3121 242
rect 3157 236 3169 242
rect 3251 236 3263 242
rect 3301 236 3313 242
rect 3363 236 3375 242
rect 3411 236 3423 242
rect 3469 236 3481 242
rect 3531 236 3543 242
rect 3571 236 3583 242
rect 3619 236 3631 242
rect 3677 236 3689 242
rect 3725 236 3737 242
rect 3787 236 3799 242
rect 3837 236 3849 242
rect 3917 236 3929 242
rect 3997 236 4009 242
rect 4037 236 4049 242
rect 1586 178 1604 180
rect 1073 104 1081 139
rect 1173 104 1181 139
rect 517 18 529 24
rect 557 18 569 24
rect 637 18 649 24
rect 771 18 783 24
rect 817 18 829 24
rect 896 18 908 24
rect 946 18 958 24
rect 1011 18 1023 24
rect 1042 18 1054 24
rect 1092 18 1104 24
rect 1298 72 1305 127
rect 1574 169 1604 178
rect 1596 141 1604 169
rect 1654 153 1662 196
rect 1869 188 1881 196
rect 1857 182 1881 188
rect 1921 190 1929 216
rect 2011 196 2021 206
rect 1921 184 1943 190
rect 1786 178 1804 180
rect 1398 72 1405 127
rect 1454 104 1462 139
rect 1774 169 1804 178
rect 1796 141 1804 169
rect 1258 66 1305 72
rect 1258 64 1269 66
rect 1142 18 1154 24
rect 1192 18 1204 24
rect 1297 64 1305 66
rect 1358 66 1405 72
rect 1358 64 1369 66
rect 1397 64 1405 66
rect 1483 98 1523 104
rect 1511 96 1523 98
rect 1598 72 1605 127
rect 1654 104 1662 139
rect 1857 133 1865 182
rect 1940 178 1943 184
rect 1558 66 1605 72
rect 1558 64 1569 66
rect 1597 64 1605 66
rect 1683 98 1723 104
rect 1711 96 1723 98
rect 1798 72 1805 127
rect 1940 122 1947 178
rect 1961 153 1969 196
rect 1967 139 1969 153
rect 1758 66 1805 72
rect 1758 64 1769 66
rect 1797 64 1805 66
rect 1857 64 1865 119
rect 1940 116 1943 122
rect 1917 110 1943 116
rect 1917 64 1925 110
rect 1961 104 1969 139
rect 2011 153 2019 196
rect 2071 186 2083 196
rect 2045 178 2083 186
rect 2101 190 2109 216
rect 2101 184 2123 190
rect 2120 178 2123 184
rect 2011 139 2013 153
rect 2011 104 2019 139
rect 2054 64 2062 178
rect 2120 122 2127 178
rect 2141 153 2149 196
rect 2409 196 2437 202
rect 2226 178 2244 180
rect 2214 169 2244 178
rect 2147 139 2149 153
rect 2236 141 2244 169
rect 2120 116 2123 122
rect 2097 110 2123 116
rect 2097 64 2105 110
rect 2141 104 2149 139
rect 2313 153 2320 196
rect 2397 193 2449 196
rect 2514 196 2540 207
rect 2609 196 2637 202
rect 2457 182 2465 196
rect 2440 175 2465 182
rect 2439 153 2447 175
rect 2514 153 2522 196
rect 2597 193 2649 196
rect 2657 182 2665 196
rect 2640 175 2665 182
rect 2639 153 2647 175
rect 2716 161 2724 216
rect 2806 178 2824 180
rect 2794 169 2824 178
rect 2238 72 2245 127
rect 2321 116 2327 139
rect 2321 110 2348 116
rect 2336 104 2348 110
rect 2433 104 2441 139
rect 2514 104 2522 139
rect 2633 104 2641 139
rect 2198 66 2245 72
rect 2198 64 2209 66
rect 2237 64 2245 66
rect 2289 96 2317 102
rect 2329 24 2357 30
rect 2543 98 2583 104
rect 2571 96 2583 98
rect 2716 64 2724 147
rect 2816 141 2824 169
rect 2876 161 2884 216
rect 2960 216 2973 222
rect 2960 210 2967 216
rect 3025 204 3032 216
rect 2818 72 2825 127
rect 2778 66 2825 72
rect 2778 64 2789 66
rect 1237 18 1249 24
rect 1277 18 1289 24
rect 1337 18 1349 24
rect 1377 18 1389 24
rect 1491 18 1503 24
rect 1537 18 1549 24
rect 1577 18 1589 24
rect 1691 18 1703 24
rect 1737 18 1749 24
rect 1777 18 1789 24
rect 1837 18 1849 24
rect 1877 18 1889 24
rect 1939 18 1951 24
rect 2027 18 2039 24
rect 2071 18 2083 24
rect 2119 18 2131 24
rect 2177 18 2189 24
rect 2217 18 2229 24
rect 2297 18 2309 24
rect 2402 18 2414 24
rect 2452 18 2464 24
rect 2551 18 2563 24
rect 2602 18 2614 24
rect 2652 18 2664 24
rect 2817 64 2825 66
rect 2876 64 2884 147
rect 2921 112 2927 196
rect 3011 197 3032 204
rect 3082 210 3089 216
rect 3082 202 3093 210
rect 2979 186 2986 192
rect 3047 186 3053 188
rect 2979 180 3053 186
rect 3135 181 3143 196
rect 2979 172 2986 180
rect 2940 164 2974 172
rect 2940 159 2946 164
rect 2966 146 2993 153
rect 2921 104 2983 112
rect 2995 108 3039 114
rect 2977 90 3015 98
rect 3033 94 3039 108
rect 3047 108 3053 180
rect 3127 167 3143 181
rect 3113 153 3127 167
rect 3047 102 3087 108
rect 3107 108 3121 116
rect 3135 104 3143 167
rect 3176 161 3184 216
rect 3236 161 3244 216
rect 3320 216 3333 222
rect 3320 210 3327 216
rect 3385 204 3392 216
rect 2977 84 2985 90
rect 3033 88 3063 94
rect 3081 84 3087 102
rect 2967 70 2985 84
rect 3013 70 3035 82
rect 2977 64 2985 70
rect 3027 64 3039 70
rect 3081 44 3093 78
rect 3176 64 3184 147
rect 3236 64 3244 147
rect 3281 112 3287 196
rect 3371 197 3392 204
rect 3442 210 3449 216
rect 3442 202 3453 210
rect 3339 186 3346 192
rect 3407 186 3413 188
rect 3339 180 3413 186
rect 3495 181 3503 196
rect 3339 172 3346 180
rect 3300 164 3334 172
rect 3300 159 3306 164
rect 3326 146 3353 153
rect 3281 104 3343 112
rect 3355 108 3399 114
rect 3337 90 3375 98
rect 3393 94 3399 108
rect 3407 108 3413 180
rect 3487 167 3503 181
rect 3473 153 3487 167
rect 3407 102 3447 108
rect 3467 108 3481 116
rect 3495 104 3503 167
rect 3553 173 3560 216
rect 3767 216 3780 222
rect 3651 210 3658 216
rect 3647 202 3658 210
rect 3708 204 3715 216
rect 3773 210 3780 216
rect 3597 181 3605 196
rect 3708 197 3729 204
rect 3687 186 3693 188
rect 3754 186 3761 192
rect 3597 167 3613 181
rect 3687 180 3761 186
rect 3553 111 3560 159
rect 3337 84 3345 90
rect 3393 88 3423 94
rect 3441 84 3447 102
rect 3327 70 3345 84
rect 3373 70 3395 82
rect 3337 64 3345 70
rect 3387 64 3399 70
rect 3441 44 3453 78
rect 3543 104 3560 111
rect 3597 104 3605 167
rect 3613 153 3627 167
rect 3619 108 3633 116
rect 3687 108 3693 180
rect 3754 172 3761 180
rect 3766 164 3800 172
rect 3794 159 3800 164
rect 3747 146 3774 153
rect 3653 102 3693 108
rect 3701 108 3745 114
rect 3653 84 3659 102
rect 3701 94 3707 108
rect 3813 112 3819 196
rect 3856 161 3864 216
rect 3909 196 3937 202
rect 3897 193 3949 196
rect 4077 236 4089 242
rect 4117 236 4129 242
rect 4171 236 4183 242
rect 4211 236 4223 242
rect 4257 236 4269 242
rect 4389 236 4401 242
rect 4451 236 4463 242
rect 3957 182 3965 196
rect 3940 175 3965 182
rect 3757 104 3819 112
rect 3677 88 3707 94
rect 3725 90 3763 98
rect 3755 84 3763 90
rect 3647 44 3659 78
rect 3705 70 3727 82
rect 3755 70 3773 84
rect 3701 64 3713 70
rect 3755 64 3763 70
rect 3856 64 3864 147
rect 3939 153 3947 175
rect 4020 173 4027 216
rect 4100 173 4107 216
rect 3933 104 3941 139
rect 4020 111 4027 159
rect 4100 111 4107 159
rect 4193 173 4200 216
rect 4249 196 4277 202
rect 4237 193 4289 196
rect 4477 236 4489 242
rect 4517 236 4529 242
rect 4559 236 4571 242
rect 4671 236 4683 242
rect 4297 182 4305 196
rect 4359 188 4371 196
rect 4359 182 4383 188
rect 4280 175 4305 182
rect 4193 111 4200 159
rect 4279 153 4287 175
rect 4020 104 4037 111
rect 4100 104 4117 111
rect 2697 18 2709 24
rect 2757 18 2769 24
rect 2797 18 2809 24
rect 2857 18 2869 24
rect 2941 18 2953 24
rect 3007 18 3019 24
rect 3053 18 3065 24
rect 3111 18 3123 24
rect 3157 18 3169 24
rect 3251 18 3263 24
rect 3301 18 3313 24
rect 3367 18 3379 24
rect 3413 18 3425 24
rect 3471 18 3483 24
rect 3571 18 3583 24
rect 3617 18 3629 24
rect 3675 18 3687 24
rect 3721 18 3733 24
rect 3787 18 3799 24
rect 3837 18 3849 24
rect 3902 18 3914 24
rect 3952 18 3964 24
rect 4183 104 4200 111
rect 4273 104 4281 139
rect 4375 133 4383 182
rect 4436 161 4444 216
rect 4500 173 4507 216
rect 4699 236 4711 242
rect 4589 188 4601 196
rect 3997 18 4009 24
rect 4077 18 4089 24
rect 4211 18 4223 24
rect 4375 64 4383 119
rect 4436 64 4444 147
rect 4500 111 4507 159
rect 4577 182 4601 188
rect 4577 133 4585 182
rect 4656 161 4664 216
rect 4729 188 4741 196
rect 4717 182 4741 188
rect 4500 104 4517 111
rect 4242 18 4254 24
rect 4292 18 4304 24
rect 4351 18 4363 24
rect 4391 18 4403 24
rect 4451 18 4463 24
rect 4577 64 4585 119
rect 4656 64 4664 147
rect 4717 133 4725 182
rect 4717 64 4725 119
rect 4477 18 4489 24
rect 4557 18 4569 24
rect 4597 18 4609 24
rect 4671 18 4683 24
rect 4697 18 4709 24
rect 4737 18 4749 24
rect -62 16 4776 18
rect -62 4 4 16
rect -62 2 4776 4
rect 4782 2 4842 242
<< m2contact >>
rect 33 4459 47 4473
rect 53 4467 67 4481
rect 73 4479 87 4493
rect 93 4467 107 4481
rect 413 4467 427 4481
rect 433 4479 447 4493
rect 453 4467 467 4481
rect 493 4493 507 4507
rect 133 4447 147 4461
rect 153 4439 167 4453
rect 193 4439 207 4453
rect 213 4439 227 4453
rect 253 4439 267 4453
rect 273 4447 287 4461
rect 333 4447 347 4461
rect 473 4459 487 4473
rect 173 4419 187 4433
rect 233 4419 247 4433
rect 353 4439 367 4453
rect 393 4439 407 4453
rect 373 4419 387 4433
rect 513 4459 527 4473
rect 533 4467 547 4481
rect 553 4459 567 4473
rect 613 4459 627 4473
rect 633 4467 647 4481
rect 653 4459 667 4473
rect 493 4433 507 4447
rect 573 4439 587 4453
rect 673 4439 687 4453
rect 733 4447 747 4461
rect 753 4439 767 4453
rect 793 4439 807 4453
rect 813 4439 827 4453
rect 853 4439 867 4453
rect 873 4447 887 4461
rect 913 4447 927 4461
rect 1093 4467 1107 4481
rect 1113 4479 1127 4493
rect 1133 4467 1147 4481
rect 773 4419 787 4433
rect 833 4419 847 4433
rect 933 4439 947 4453
rect 953 4447 967 4461
rect 993 4439 1007 4453
rect 1033 4439 1047 4453
rect 1053 4447 1067 4461
rect 1153 4459 1167 4473
rect 1013 4419 1027 4433
rect 1213 4447 1227 4461
rect 1313 4479 1327 4493
rect 1233 4439 1247 4453
rect 1253 4447 1267 4461
rect 1293 4459 1307 4473
rect 1333 4459 1347 4473
rect 1393 4459 1407 4473
rect 1413 4467 1427 4481
rect 1433 4459 1447 4473
rect 1373 4439 1387 4453
rect 1473 4447 1487 4461
rect 1553 4479 1567 4493
rect 1493 4439 1507 4453
rect 1513 4447 1527 4461
rect 1533 4459 1547 4473
rect 1573 4459 1587 4473
rect 1613 4439 1627 4453
rect 1653 4439 1667 4453
rect 1673 4447 1687 4461
rect 1733 4459 1747 4473
rect 1753 4467 1767 4481
rect 1773 4479 1787 4493
rect 1793 4467 1807 4481
rect 1813 4479 1827 4493
rect 1833 4467 1847 4481
rect 1893 4467 1907 4481
rect 1913 4479 1927 4493
rect 1933 4467 1947 4481
rect 1953 4479 1967 4493
rect 1973 4467 1987 4481
rect 2053 4479 2067 4493
rect 2113 4479 2127 4493
rect 2753 4516 2767 4530
rect 1633 4419 1647 4433
rect 1993 4459 2007 4473
rect 2033 4459 2047 4473
rect 2073 4459 2087 4473
rect 2133 4467 2147 4481
rect 2173 4459 2187 4473
rect 2193 4467 2207 4481
rect 2213 4459 2227 4473
rect 2293 4459 2307 4473
rect 2313 4467 2327 4481
rect 2333 4459 2347 4473
rect 2353 4467 2367 4481
rect 2393 4479 2407 4493
rect 2373 4459 2387 4473
rect 2413 4459 2427 4473
rect 2233 4439 2247 4453
rect 2453 4467 2467 4481
rect 2493 4467 2507 4481
rect 2513 4479 2527 4493
rect 2533 4467 2547 4481
rect 2553 4459 2567 4473
rect 2613 4459 2627 4473
rect 2633 4467 2647 4481
rect 2653 4459 2667 4473
rect 2673 4467 2687 4481
rect 2693 4459 2707 4473
rect 2893 4516 2907 4530
rect 2793 4459 2807 4473
rect 2833 4459 2847 4473
rect 2913 4487 2927 4501
rect 2893 4422 2907 4436
rect 2973 4467 2987 4481
rect 2993 4479 3007 4493
rect 2753 4390 2767 4404
rect 2893 4384 2907 4398
rect 3053 4459 3067 4473
rect 3073 4467 3087 4481
rect 3093 4459 3107 4473
rect 3033 4439 3047 4453
rect 3133 4513 3147 4527
rect 3153 4479 3167 4493
rect 3133 4459 3147 4473
rect 3113 4433 3127 4447
rect 3173 4459 3187 4473
rect 3233 4459 3247 4473
rect 3253 4467 3267 4481
rect 3333 4479 3347 4493
rect 3473 4516 3487 4530
rect 3613 4516 3627 4530
rect 3273 4459 3287 4473
rect 3313 4459 3327 4473
rect 3213 4439 3227 4453
rect 3353 4459 3367 4473
rect 3393 4467 3407 4481
rect 3413 4479 3427 4493
rect 3453 4487 3467 4501
rect 3473 4422 3487 4436
rect 3533 4459 3547 4473
rect 3573 4459 3587 4473
rect 3673 4459 3687 4473
rect 3693 4467 3707 4481
rect 3713 4459 3727 4473
rect 3733 4439 3747 4453
rect 3773 4447 3787 4461
rect 3873 4467 3887 4481
rect 3793 4439 3807 4453
rect 3813 4447 3827 4461
rect 3473 4384 3487 4398
rect 3613 4390 3627 4404
rect 4013 4467 4027 4481
rect 4073 4459 4087 4473
rect 4113 4459 4127 4473
rect 4133 4447 4147 4461
rect 4213 4479 4227 4493
rect 4413 4516 4427 4530
rect 4553 4516 4567 4530
rect 4233 4467 4247 4481
rect 4153 4439 4167 4453
rect 4173 4447 4187 4461
rect 4273 4459 4287 4473
rect 4293 4467 4307 4481
rect 4313 4459 4327 4473
rect 4393 4487 4407 4501
rect 4333 4439 4347 4453
rect 4413 4422 4427 4436
rect 4473 4459 4487 4473
rect 4513 4459 4527 4473
rect 4613 4459 4627 4473
rect 4653 4459 4667 4473
rect 4413 4384 4427 4398
rect 4553 4390 4567 4404
rect 4693 4447 4707 4461
rect 4713 4439 4727 4453
rect 4733 4447 4747 4461
rect 33 4199 47 4213
rect 53 4207 67 4221
rect 73 4199 87 4213
rect 93 4179 107 4193
rect 113 4167 127 4181
rect 133 4179 147 4193
rect 153 4187 167 4201
rect 213 4199 227 4213
rect 233 4207 247 4221
rect 253 4199 267 4213
rect 293 4187 307 4201
rect 373 4207 387 4221
rect 513 4207 527 4221
rect 333 4187 347 4201
rect 393 4187 407 4201
rect 313 4167 327 4181
rect 413 4179 427 4193
rect 433 4187 447 4201
rect 453 4187 467 4201
rect 473 4179 487 4193
rect 493 4187 507 4201
rect 573 4179 587 4193
rect 633 4187 647 4201
rect 793 4227 807 4241
rect 773 4207 787 4221
rect 813 4207 827 4221
rect 833 4199 847 4213
rect 1053 4227 1067 4241
rect 1113 4227 1127 4241
rect 593 4167 607 4181
rect 653 4179 667 4193
rect 673 4167 687 4181
rect 693 4179 707 4193
rect 733 4179 747 4193
rect 753 4167 767 4181
rect 893 4187 907 4201
rect 913 4179 927 4193
rect 933 4187 947 4201
rect 953 4179 967 4193
rect 973 4187 987 4201
rect 1013 4199 1027 4213
rect 1033 4207 1047 4221
rect 1073 4207 1087 4221
rect 1093 4207 1107 4221
rect 1133 4207 1147 4221
rect 1153 4199 1167 4213
rect 1213 4199 1227 4213
rect 1233 4207 1247 4221
rect 1333 4227 1347 4241
rect 1473 4227 1487 4241
rect 1253 4199 1267 4213
rect 1293 4199 1307 4213
rect 1313 4207 1327 4221
rect 1353 4207 1367 4221
rect 1393 4199 1407 4213
rect 1413 4207 1427 4221
rect 1433 4199 1447 4213
rect 1453 4207 1467 4221
rect 1493 4207 1507 4221
rect 1513 4199 1527 4213
rect 1573 4187 1587 4201
rect 1613 4187 1627 4201
rect 1653 4187 1667 4201
rect 1773 4207 1787 4221
rect 1693 4187 1707 4201
rect 1713 4187 1727 4201
rect 1593 4167 1607 4181
rect 1673 4167 1687 4181
rect 1733 4179 1747 4193
rect 1753 4187 1767 4201
rect 1833 4199 1847 4213
rect 1853 4207 1867 4221
rect 1873 4199 1887 4213
rect 1973 4227 1987 4241
rect 1953 4207 1967 4221
rect 1993 4207 2007 4221
rect 2073 4227 2087 4241
rect 2013 4199 2027 4213
rect 2053 4207 2067 4221
rect 2093 4207 2107 4221
rect 2193 4256 2207 4270
rect 2333 4262 2347 4276
rect 2113 4199 2127 4213
rect 1893 4167 1907 4181
rect 1913 4179 1927 4193
rect 2233 4187 2247 4201
rect 2273 4187 2287 4201
rect 2333 4224 2347 4238
rect 2393 4187 2407 4201
rect 2353 4159 2367 4173
rect 2193 4130 2207 4144
rect 2433 4187 2447 4201
rect 2653 4262 2667 4276
rect 2793 4256 2807 4270
rect 2333 4130 2347 4144
rect 2493 4179 2507 4193
rect 2553 4187 2567 4201
rect 2593 4187 2607 4201
rect 2513 4167 2527 4181
rect 2573 4167 2587 4181
rect 2653 4224 2667 4238
rect 2633 4159 2647 4173
rect 2713 4187 2727 4201
rect 2753 4187 2767 4201
rect 2653 4130 2667 4144
rect 2853 4167 2867 4181
rect 2873 4179 2887 4193
rect 2933 4187 2947 4201
rect 3453 4256 3467 4270
rect 3593 4262 3607 4276
rect 3053 4207 3067 4221
rect 2973 4187 2987 4201
rect 2993 4187 3007 4201
rect 2793 4130 2807 4144
rect 2953 4167 2967 4181
rect 3013 4179 3027 4193
rect 3033 4187 3047 4201
rect 3093 4199 3107 4213
rect 3113 4207 3127 4221
rect 3133 4199 3147 4213
rect 3193 4199 3207 4213
rect 3213 4207 3227 4221
rect 3233 4199 3247 4213
rect 3273 4199 3287 4213
rect 3293 4207 3307 4221
rect 3313 4199 3327 4213
rect 3333 4187 3347 4201
rect 3373 4187 3387 4201
rect 3353 4167 3367 4181
rect 3493 4187 3507 4201
rect 3533 4187 3547 4201
rect 3593 4224 3607 4238
rect 3853 4262 3867 4276
rect 3993 4256 4007 4270
rect 3673 4199 3687 4213
rect 3693 4207 3707 4221
rect 3613 4159 3627 4173
rect 3453 4130 3467 4144
rect 3713 4199 3727 4213
rect 3733 4187 3747 4201
rect 3773 4187 3787 4201
rect 3753 4167 3767 4181
rect 3593 4130 3607 4144
rect 3853 4224 3867 4238
rect 3833 4159 3847 4173
rect 3913 4187 3927 4201
rect 3953 4187 3967 4201
rect 3853 4130 3867 4144
rect 4053 4187 4067 4201
rect 4533 4262 4547 4276
rect 4673 4256 4687 4270
rect 4093 4187 4107 4201
rect 4153 4187 4167 4201
rect 4073 4167 4087 4181
rect 3993 4130 4007 4144
rect 4173 4179 4187 4193
rect 4193 4167 4207 4181
rect 4213 4179 4227 4193
rect 4233 4187 4247 4201
rect 4273 4187 4287 4201
rect 4333 4187 4347 4201
rect 4373 4187 4387 4201
rect 4413 4187 4427 4201
rect 4353 4167 4367 4181
rect 4433 4179 4447 4193
rect 4453 4167 4467 4181
rect 4473 4179 4487 4193
rect 4533 4224 4547 4238
rect 4513 4159 4527 4173
rect 4593 4187 4607 4201
rect 4633 4187 4647 4201
rect 4533 4130 4547 4144
rect 4673 4130 4687 4144
rect 33 3967 47 3981
rect 53 3959 67 3973
rect 73 3967 87 3981
rect 93 3967 107 3981
rect 113 3959 127 3973
rect 133 3967 147 3981
rect 193 3967 207 3981
rect 213 3959 227 3973
rect 233 3967 247 3981
rect 293 3979 307 3993
rect 313 3987 327 4001
rect 333 3979 347 3993
rect 353 3987 367 4001
rect 373 3999 387 4013
rect 393 3987 407 4001
rect 493 3999 507 4013
rect 413 3979 427 3993
rect 473 3979 487 3993
rect 273 3959 287 3973
rect 513 3979 527 3993
rect 533 3967 547 3981
rect 553 3959 567 3973
rect 573 3967 587 3981
rect 613 3979 627 3993
rect 633 3987 647 4001
rect 653 3979 667 3993
rect 673 3959 687 3973
rect 733 3967 747 3981
rect 753 3959 767 3973
rect 793 3959 807 3973
rect 813 3959 827 3973
rect 853 3959 867 3973
rect 873 3967 887 3981
rect 953 3979 967 3993
rect 973 3987 987 4001
rect 993 3979 1007 3993
rect 1013 3979 1027 3993
rect 1033 3987 1047 4001
rect 1053 3979 1067 3993
rect 1133 3987 1147 4001
rect 1153 3999 1167 4013
rect 773 3939 787 3953
rect 833 3939 847 3953
rect 933 3959 947 3973
rect 1073 3959 1087 3973
rect 1273 3999 1287 4013
rect 1293 3987 1307 4001
rect 1193 3967 1207 3981
rect 1213 3959 1227 3973
rect 1253 3959 1267 3973
rect 1233 3939 1247 3953
rect 1333 3959 1347 3973
rect 1373 3959 1387 3973
rect 1393 3967 1407 3981
rect 1353 3939 1367 3953
rect 1433 3959 1447 3973
rect 1473 3959 1487 3973
rect 1493 3967 1507 3981
rect 1533 3967 1547 3981
rect 1653 3999 1667 4013
rect 1453 3939 1467 3953
rect 1553 3959 1567 3973
rect 1573 3967 1587 3981
rect 1633 3979 1647 3993
rect 1673 3979 1687 3993
rect 1713 3979 1727 3993
rect 1733 3967 1747 3981
rect 1773 3979 1787 3993
rect 1833 3979 1847 3993
rect 1853 3987 1867 4001
rect 1913 3999 1927 4013
rect 1873 3979 1887 3993
rect 1893 3979 1907 3993
rect 1813 3959 1827 3973
rect 1933 3979 1947 3993
rect 1993 3987 2007 4001
rect 2013 3999 2027 4013
rect 2033 3979 2047 3993
rect 2053 3987 2067 4001
rect 2133 3999 2147 4013
rect 2073 3979 2087 3993
rect 2153 3987 2167 4001
rect 2093 3959 2107 3973
rect 2193 3967 2207 3981
rect 2693 4036 2707 4050
rect 2213 3959 2227 3973
rect 2233 3967 2247 3981
rect 2273 3959 2287 3973
rect 2313 3959 2327 3973
rect 2333 3967 2347 3981
rect 2373 3979 2387 3993
rect 2293 3939 2307 3953
rect 2413 3979 2427 3993
rect 2473 3987 2487 4001
rect 2613 3987 2627 4001
rect 2833 4036 2847 4050
rect 2733 3979 2747 3993
rect 2773 3979 2787 3993
rect 2853 4007 2867 4021
rect 2833 3942 2847 3956
rect 2893 3999 2907 4013
rect 2913 3987 2927 4001
rect 2693 3910 2707 3924
rect 2833 3904 2847 3918
rect 2953 3979 2967 3993
rect 2973 3987 2987 4001
rect 3073 3999 3087 4013
rect 2993 3979 3007 3993
rect 3053 3979 3067 3993
rect 3013 3959 3027 3973
rect 3093 3979 3107 3993
rect 3133 3967 3147 3981
rect 3153 3959 3167 3973
rect 3173 3967 3187 3981
rect 3233 3979 3247 3993
rect 3253 3987 3267 4001
rect 3273 3999 3287 4013
rect 3293 3987 3307 4001
rect 3313 3979 3327 3993
rect 3453 3999 3467 4013
rect 3593 4036 3607 4050
rect 3733 4036 3747 4050
rect 3353 3967 3367 3981
rect 3373 3979 3387 3993
rect 3433 3979 3447 3993
rect 3473 3979 3487 3993
rect 3513 3987 3527 4001
rect 3533 3999 3547 4013
rect 3573 4007 3587 4021
rect 3593 3942 3607 3956
rect 3653 3979 3667 3993
rect 3693 3979 3707 3993
rect 3813 3979 3827 3993
rect 3833 3987 3847 4001
rect 3853 3999 3867 4013
rect 3873 3987 3887 4001
rect 3913 3999 3927 4013
rect 3893 3979 3907 3993
rect 4013 3999 4027 4013
rect 3933 3979 3947 3993
rect 3993 3979 4007 3993
rect 4033 3979 4047 3993
rect 4053 3979 4067 3993
rect 3593 3904 3607 3918
rect 3733 3910 3747 3924
rect 4093 3967 4107 3981
rect 4113 3979 4127 3993
rect 4153 3979 4167 3993
rect 4173 3987 4187 4001
rect 4193 3979 4207 3993
rect 4333 4013 4347 4027
rect 4293 3979 4307 3993
rect 4313 3987 4327 4001
rect 4333 3979 4347 3993
rect 4213 3959 4227 3973
rect 4273 3959 4287 3973
rect 4453 4036 4467 4050
rect 4593 4036 4607 4050
rect 4373 3987 4387 4001
rect 4393 3999 4407 4013
rect 4433 4007 4447 4021
rect 4353 3953 4367 3967
rect 4453 3942 4467 3956
rect 4513 3979 4527 3993
rect 4553 3979 4567 3993
rect 4653 3999 4667 4013
rect 4673 3987 4687 4001
rect 4453 3904 4467 3918
rect 4593 3910 4607 3924
rect 33 3707 47 3721
rect 153 3727 167 3741
rect 73 3707 87 3721
rect 93 3707 107 3721
rect 53 3687 67 3701
rect 113 3699 127 3713
rect 133 3707 147 3721
rect 213 3699 227 3713
rect 273 3707 287 3721
rect 233 3687 247 3701
rect 293 3699 307 3713
rect 313 3687 327 3701
rect 333 3699 347 3713
rect 373 3707 387 3721
rect 393 3719 407 3733
rect 433 3707 447 3721
rect 473 3719 487 3733
rect 493 3727 507 3741
rect 513 3719 527 3733
rect 553 3753 567 3767
rect 553 3719 567 3733
rect 573 3727 587 3741
rect 533 3673 547 3687
rect 593 3719 607 3733
rect 753 3753 767 3767
rect 733 3727 747 3741
rect 613 3687 627 3701
rect 633 3699 647 3713
rect 673 3707 687 3721
rect 693 3699 707 3713
rect 713 3707 727 3721
rect 733 3693 747 3707
rect 773 3719 787 3733
rect 793 3727 807 3741
rect 913 3747 927 3761
rect 813 3719 827 3733
rect 873 3719 887 3733
rect 893 3727 907 3741
rect 933 3727 947 3741
rect 1073 3747 1087 3761
rect 1053 3727 1067 3741
rect 1093 3727 1107 3741
rect 953 3699 967 3713
rect 973 3687 987 3701
rect 993 3699 1007 3713
rect 1013 3707 1027 3721
rect 1113 3719 1127 3733
rect 1153 3699 1167 3713
rect 1173 3687 1187 3701
rect 1193 3699 1207 3713
rect 1213 3707 1227 3721
rect 1373 3747 1387 3761
rect 1333 3719 1347 3733
rect 1353 3727 1367 3741
rect 1393 3727 1407 3741
rect 1253 3687 1267 3701
rect 1273 3699 1287 3713
rect 1493 3727 1507 3741
rect 1433 3699 1447 3713
rect 1513 3707 1527 3721
rect 1453 3687 1467 3701
rect 1533 3699 1547 3713
rect 1553 3707 1567 3721
rect 1593 3699 1607 3713
rect 1613 3687 1627 3701
rect 1633 3699 1647 3713
rect 1653 3687 1667 3701
rect 1673 3699 1687 3713
rect 1693 3707 1707 3721
rect 1733 3707 1747 3721
rect 1773 3707 1787 3721
rect 1833 3707 1847 3721
rect 1933 3719 1947 3733
rect 1953 3727 1967 3741
rect 1753 3687 1767 3701
rect 1853 3699 1867 3713
rect 1873 3687 1887 3701
rect 1893 3699 1907 3713
rect 1973 3719 1987 3733
rect 2013 3707 2027 3721
rect 1993 3687 2007 3701
rect 2413 3776 2427 3790
rect 2553 3782 2567 3796
rect 2053 3699 2067 3713
rect 2093 3707 2107 3721
rect 2133 3707 2147 3721
rect 2193 3699 2207 3713
rect 2333 3699 2347 3713
rect 2453 3707 2467 3721
rect 2493 3707 2507 3721
rect 2553 3744 2567 3758
rect 2633 3727 2647 3741
rect 2573 3679 2587 3693
rect 2653 3707 2667 3721
rect 2673 3699 2687 3713
rect 2693 3707 2707 3721
rect 2733 3699 2747 3713
rect 2793 3707 2807 3721
rect 2833 3707 2847 3721
rect 2873 3707 2887 3721
rect 2913 3707 2927 3721
rect 2953 3707 2967 3721
rect 2993 3707 3007 3721
rect 3193 3727 3207 3741
rect 2413 3650 2427 3664
rect 2553 3650 2567 3664
rect 2753 3687 2767 3701
rect 2813 3687 2827 3701
rect 2893 3687 2907 3701
rect 2973 3687 2987 3701
rect 3013 3687 3027 3701
rect 3033 3699 3047 3713
rect 3093 3699 3107 3713
rect 3133 3707 3147 3721
rect 3113 3687 3127 3701
rect 3153 3699 3167 3713
rect 3173 3707 3187 3721
rect 3253 3707 3267 3721
rect 3273 3699 3287 3713
rect 3293 3687 3307 3701
rect 3313 3699 3327 3713
rect 3333 3699 3347 3713
rect 3353 3687 3367 3701
rect 3373 3699 3387 3713
rect 3393 3707 3407 3721
rect 3433 3687 3447 3701
rect 3453 3699 3467 3713
rect 3493 3707 3507 3721
rect 3833 3776 3847 3790
rect 3973 3782 3987 3796
rect 3533 3719 3547 3733
rect 3653 3727 3667 3741
rect 3753 3727 3767 3741
rect 3553 3707 3567 3721
rect 3593 3707 3607 3721
rect 3613 3699 3627 3713
rect 3633 3707 3647 3721
rect 3693 3707 3707 3721
rect 3713 3699 3727 3713
rect 3733 3707 3747 3721
rect 3873 3707 3887 3721
rect 3913 3707 3927 3721
rect 3973 3744 3987 3758
rect 4333 3782 4347 3796
rect 4473 3776 4487 3790
rect 4033 3707 4047 3721
rect 3993 3679 4007 3693
rect 3833 3650 3847 3664
rect 4073 3707 4087 3721
rect 4133 3707 4147 3721
rect 3973 3650 3987 3664
rect 4173 3707 4187 3721
rect 4153 3687 4167 3701
rect 4193 3699 4207 3713
rect 4213 3687 4227 3701
rect 4233 3699 4247 3713
rect 4253 3707 4267 3721
rect 4333 3744 4347 3758
rect 4313 3679 4327 3693
rect 4393 3707 4407 3721
rect 4433 3707 4447 3721
rect 4333 3650 4347 3664
rect 4533 3707 4547 3721
rect 4573 3707 4587 3721
rect 4473 3650 4487 3664
rect 4633 3699 4647 3713
rect 4653 3687 4667 3701
rect 4673 3687 4687 3701
rect 4693 3699 4707 3713
rect 133 3556 147 3570
rect 33 3487 47 3501
rect 53 3479 67 3493
rect 73 3487 87 3501
rect 273 3556 287 3570
rect 173 3499 187 3513
rect 213 3499 227 3513
rect 293 3527 307 3541
rect 273 3462 287 3476
rect 353 3507 367 3521
rect 373 3519 387 3533
rect 133 3430 147 3444
rect 273 3424 287 3438
rect 413 3487 427 3501
rect 433 3479 447 3493
rect 453 3487 467 3501
rect 513 3499 527 3513
rect 533 3507 547 3521
rect 553 3499 567 3513
rect 613 3499 627 3513
rect 633 3507 647 3521
rect 653 3499 667 3513
rect 493 3479 507 3493
rect 593 3479 607 3493
rect 673 3487 687 3501
rect 693 3479 707 3493
rect 713 3487 727 3501
rect 753 3499 767 3513
rect 773 3507 787 3521
rect 793 3499 807 3513
rect 813 3507 827 3521
rect 873 3519 887 3533
rect 833 3499 847 3513
rect 893 3507 907 3521
rect 953 3553 967 3567
rect 1033 3507 1047 3521
rect 1053 3519 1067 3533
rect 1073 3507 1087 3521
rect 1513 3556 1527 3570
rect 1153 3519 1167 3533
rect 953 3487 967 3501
rect 1093 3499 1107 3513
rect 1133 3499 1147 3513
rect 933 3453 947 3467
rect 973 3479 987 3493
rect 1013 3479 1027 3493
rect 993 3459 1007 3473
rect 1173 3499 1187 3513
rect 1213 3487 1227 3501
rect 1233 3479 1247 3493
rect 1253 3487 1267 3501
rect 1293 3487 1307 3501
rect 1313 3479 1327 3493
rect 1333 3487 1347 3501
rect 1373 3499 1387 3513
rect 1393 3507 1407 3521
rect 1413 3499 1427 3513
rect 1433 3479 1447 3493
rect 1653 3556 1667 3570
rect 1553 3499 1567 3513
rect 1593 3499 1607 3513
rect 1673 3527 1687 3541
rect 1653 3462 1667 3476
rect 1733 3487 1747 3501
rect 1753 3479 1767 3493
rect 1773 3487 1787 3501
rect 1793 3499 1807 3513
rect 1813 3507 1827 3521
rect 1833 3499 1847 3513
rect 1893 3507 1907 3521
rect 1913 3499 1927 3513
rect 1513 3430 1527 3444
rect 1653 3424 1667 3438
rect 1853 3479 1867 3493
rect 1973 3487 1987 3501
rect 1993 3479 2007 3493
rect 2013 3487 2027 3501
rect 2053 3499 2067 3513
rect 2073 3487 2087 3501
rect 2113 3499 2127 3513
rect 2133 3487 2147 3501
rect 2313 3519 2327 3533
rect 2333 3507 2347 3521
rect 2373 3519 2387 3533
rect 2473 3556 2487 3570
rect 2613 3556 2627 3570
rect 2453 3527 2467 3541
rect 2393 3507 2407 3521
rect 2153 3479 2167 3493
rect 2173 3487 2187 3501
rect 2213 3479 2227 3493
rect 2253 3479 2267 3493
rect 2273 3487 2287 3501
rect 2233 3459 2247 3473
rect 2473 3462 2487 3476
rect 2533 3499 2547 3513
rect 2573 3499 2587 3513
rect 2673 3499 2687 3513
rect 2693 3507 2707 3521
rect 2713 3499 2727 3513
rect 2773 3499 2787 3513
rect 2733 3479 2747 3493
rect 2973 3556 2987 3570
rect 2813 3499 2827 3513
rect 2473 3424 2487 3438
rect 2613 3430 2627 3444
rect 2853 3487 2867 3501
rect 3113 3556 3127 3570
rect 2953 3527 2967 3541
rect 2873 3479 2887 3493
rect 2893 3487 2907 3501
rect 2973 3462 2987 3476
rect 3033 3499 3047 3513
rect 3073 3499 3087 3513
rect 3393 3533 3407 3547
rect 3213 3499 3227 3513
rect 3233 3507 3247 3521
rect 3253 3499 3267 3513
rect 3293 3507 3307 3521
rect 3313 3519 3327 3533
rect 3353 3519 3367 3533
rect 3193 3479 3207 3493
rect 2973 3424 2987 3438
rect 3113 3430 3127 3444
rect 3333 3499 3347 3513
rect 3373 3499 3387 3513
rect 3413 3519 3427 3533
rect 3433 3507 3447 3521
rect 3513 3519 3527 3533
rect 3413 3473 3427 3487
rect 3493 3499 3507 3513
rect 3533 3499 3547 3513
rect 3553 3507 3567 3521
rect 3573 3519 3587 3533
rect 3593 3507 3607 3521
rect 3993 3556 4007 3570
rect 3653 3519 3667 3533
rect 3613 3499 3627 3513
rect 3673 3499 3687 3513
rect 3713 3507 3727 3521
rect 3773 3499 3787 3513
rect 3793 3507 3807 3521
rect 3813 3499 3827 3513
rect 3833 3507 3847 3521
rect 3853 3499 3867 3513
rect 3893 3487 3907 3501
rect 4133 3556 4147 3570
rect 3973 3527 3987 3541
rect 3913 3479 3927 3493
rect 3933 3487 3947 3501
rect 3993 3462 4007 3476
rect 4053 3499 4067 3513
rect 4093 3499 4107 3513
rect 3993 3424 4007 3438
rect 4133 3430 4147 3444
rect 4233 3556 4247 3570
rect 4373 3556 4387 3570
rect 4213 3527 4227 3541
rect 4233 3462 4247 3476
rect 4293 3499 4307 3513
rect 4333 3499 4347 3513
rect 4453 3507 4467 3521
rect 4593 3507 4607 3521
rect 4633 3499 4647 3513
rect 4653 3507 4667 3521
rect 4673 3499 4687 3513
rect 4693 3479 4707 3493
rect 4233 3424 4247 3438
rect 4373 3430 4387 3444
rect 53 3296 67 3310
rect 193 3302 207 3316
rect 93 3227 107 3241
rect 133 3227 147 3241
rect 193 3264 207 3278
rect 393 3293 407 3307
rect 273 3227 287 3241
rect 293 3219 307 3233
rect 313 3227 327 3241
rect 213 3199 227 3213
rect 53 3170 67 3184
rect 333 3219 347 3233
rect 353 3227 367 3241
rect 493 3302 507 3316
rect 633 3296 647 3310
rect 393 3239 407 3253
rect 413 3247 427 3261
rect 373 3213 387 3227
rect 433 3239 447 3253
rect 493 3264 507 3278
rect 473 3199 487 3213
rect 553 3227 567 3241
rect 593 3227 607 3241
rect 193 3170 207 3184
rect 493 3170 507 3184
rect 713 3247 727 3261
rect 733 3227 747 3241
rect 753 3219 767 3233
rect 773 3227 787 3241
rect 813 3227 827 3241
rect 833 3219 847 3233
rect 853 3227 867 3241
rect 633 3170 647 3184
rect 873 3219 887 3233
rect 893 3227 907 3241
rect 913 3239 927 3253
rect 933 3247 947 3261
rect 1053 3267 1067 3281
rect 953 3239 967 3253
rect 1013 3239 1027 3253
rect 1033 3247 1047 3261
rect 1073 3247 1087 3261
rect 1113 3227 1127 3241
rect 1133 3239 1147 3253
rect 1213 3267 1227 3281
rect 1193 3247 1207 3261
rect 1233 3247 1247 3261
rect 1173 3227 1187 3241
rect 1253 3239 1267 3253
rect 1353 3247 1367 3261
rect 1293 3227 1307 3241
rect 1313 3219 1327 3233
rect 1333 3227 1347 3241
rect 1393 3239 1407 3253
rect 1413 3247 1427 3261
rect 1433 3239 1447 3253
rect 1493 3219 1507 3233
rect 1533 3227 1547 3241
rect 1553 3207 1567 3221
rect 1553 3173 1567 3187
rect 1593 3273 1607 3287
rect 1713 3293 1727 3307
rect 1773 3293 1787 3307
rect 1593 3239 1607 3253
rect 1613 3247 1627 3261
rect 1633 3239 1647 3253
rect 1713 3247 1727 3261
rect 1773 3247 1787 3261
rect 1893 3273 1907 3287
rect 1653 3227 1667 3241
rect 1673 3219 1687 3233
rect 1693 3227 1707 3241
rect 1793 3227 1807 3241
rect 1813 3219 1827 3233
rect 1833 3227 1847 3241
rect 1853 3239 1867 3253
rect 1873 3247 1887 3261
rect 1893 3239 1907 3253
rect 1993 3247 2007 3261
rect 2053 3247 2067 3261
rect 1933 3227 1947 3241
rect 1953 3219 1967 3233
rect 1973 3227 1987 3241
rect 1933 3193 1947 3207
rect 2073 3227 2087 3241
rect 2093 3219 2107 3233
rect 2113 3227 2127 3241
rect 2253 3247 2267 3261
rect 2133 3207 2147 3221
rect 2153 3219 2167 3233
rect 2193 3227 2207 3241
rect 2213 3219 2227 3233
rect 2233 3227 2247 3241
rect 2473 3302 2487 3316
rect 2613 3296 2627 3310
rect 2353 3239 2367 3253
rect 2373 3247 2387 3261
rect 2313 3219 2327 3233
rect 2333 3207 2347 3221
rect 2393 3239 2407 3253
rect 2473 3264 2487 3278
rect 2453 3199 2467 3213
rect 2533 3227 2547 3241
rect 2573 3227 2587 3241
rect 2473 3170 2487 3184
rect 2793 3302 2807 3316
rect 2933 3296 2947 3310
rect 2673 3227 2687 3241
rect 2713 3227 2727 3241
rect 2613 3170 2627 3184
rect 2793 3264 2807 3278
rect 2773 3199 2787 3213
rect 2853 3227 2867 3241
rect 2893 3227 2907 3241
rect 2793 3170 2807 3184
rect 3013 3247 3027 3261
rect 3113 3247 3127 3261
rect 3253 3247 3267 3261
rect 3313 3247 3327 3261
rect 3453 3247 3467 3261
rect 3033 3227 3047 3241
rect 3053 3219 3067 3233
rect 3073 3227 3087 3241
rect 3133 3227 3147 3241
rect 3153 3219 3167 3233
rect 3173 3227 3187 3241
rect 3193 3227 3207 3241
rect 3213 3219 3227 3233
rect 3233 3227 3247 3241
rect 3333 3227 3347 3241
rect 3353 3219 3367 3233
rect 3373 3227 3387 3241
rect 3393 3227 3407 3241
rect 3413 3219 3427 3233
rect 3433 3227 3447 3241
rect 3493 3239 3507 3253
rect 3513 3247 3527 3261
rect 2933 3170 2947 3184
rect 3533 3239 3547 3253
rect 3573 3239 3587 3253
rect 3593 3247 3607 3261
rect 3613 3239 3627 3253
rect 3653 3239 3667 3253
rect 3673 3247 3687 3261
rect 3693 3239 3707 3253
rect 3733 3239 3747 3253
rect 3753 3247 3767 3261
rect 3773 3239 3787 3253
rect 3813 3227 3827 3241
rect 3853 3227 3867 3241
rect 3913 3239 3927 3253
rect 3933 3247 3947 3261
rect 3953 3239 3967 3253
rect 3993 3227 4007 3241
rect 4033 3227 4047 3241
rect 4053 3227 4067 3241
rect 4013 3207 4027 3221
rect 4093 3227 4107 3241
rect 4213 3247 4227 3261
rect 4153 3219 4167 3233
rect 4233 3227 4247 3241
rect 4173 3207 4187 3221
rect 4253 3219 4267 3233
rect 4273 3227 4287 3241
rect 4573 3296 4587 3310
rect 4713 3302 4727 3316
rect 4413 3247 4427 3261
rect 4313 3219 4327 3233
rect 4353 3227 4367 3241
rect 4333 3207 4347 3221
rect 4373 3219 4387 3233
rect 4393 3227 4407 3241
rect 4473 3239 4487 3253
rect 4493 3247 4507 3261
rect 4513 3239 4527 3253
rect 4613 3227 4627 3241
rect 4653 3227 4667 3241
rect 4713 3264 4727 3278
rect 4733 3199 4747 3213
rect 4573 3170 4587 3184
rect 4713 3170 4727 3184
rect 33 3019 47 3033
rect 53 3027 67 3041
rect 73 3019 87 3033
rect 93 3027 107 3041
rect 273 3076 287 3090
rect 413 3076 427 3090
rect 113 3019 127 3033
rect 153 3019 167 3033
rect 173 3007 187 3021
rect 253 3047 267 3061
rect 213 3019 227 3033
rect 273 2982 287 2996
rect 333 3019 347 3033
rect 373 3019 387 3033
rect 473 3019 487 3033
rect 493 3027 507 3041
rect 513 3019 527 3033
rect 533 2999 547 3013
rect 273 2944 287 2958
rect 413 2950 427 2964
rect 533 2953 547 2967
rect 573 3053 587 3067
rect 573 3007 587 3021
rect 593 2999 607 3013
rect 613 3007 627 3021
rect 673 3007 687 3021
rect 773 3039 787 3053
rect 693 2999 707 3013
rect 713 3007 727 3021
rect 753 3019 767 3033
rect 793 3019 807 3033
rect 813 3007 827 3021
rect 833 2999 847 3013
rect 853 3007 867 3021
rect 933 3019 947 3033
rect 953 3027 967 3041
rect 973 3019 987 3033
rect 1033 3019 1047 3033
rect 1053 3027 1067 3041
rect 1133 3039 1147 3053
rect 1073 3019 1087 3033
rect 1113 3019 1127 3033
rect 913 2999 927 3013
rect 1013 2999 1027 3013
rect 1153 3019 1167 3033
rect 1213 3019 1227 3033
rect 1233 3027 1247 3041
rect 1253 3019 1267 3033
rect 1193 2999 1207 3013
rect 1273 3007 1287 3021
rect 1293 2999 1307 3013
rect 1313 3007 1327 3021
rect 1373 3019 1387 3033
rect 1393 3027 1407 3041
rect 1413 3007 1427 3021
rect 1433 2999 1447 3013
rect 1453 3007 1467 3021
rect 1493 3007 1507 3021
rect 1513 2999 1527 3013
rect 1533 3007 1547 3021
rect 1573 3019 1587 3033
rect 1613 3019 1627 3033
rect 1653 3019 1667 3033
rect 1673 3027 1687 3041
rect 1693 3019 1707 3033
rect 1753 3019 1767 3033
rect 1773 3027 1787 3041
rect 1813 3033 1827 3047
rect 1873 3039 1887 3053
rect 1793 3019 1807 3033
rect 1713 2999 1727 3013
rect 1813 2999 1827 3013
rect 1853 3019 1867 3033
rect 1893 3019 1907 3033
rect 1933 3027 1947 3041
rect 1953 3039 1967 3053
rect 1973 3027 1987 3041
rect 2033 3039 2047 3053
rect 1993 3019 2007 3033
rect 2053 3027 2067 3041
rect 1833 2973 1847 2987
rect 2093 3019 2107 3033
rect 2113 3027 2127 3041
rect 2213 3039 2227 3053
rect 2133 3019 2147 3033
rect 2193 3019 2207 3033
rect 2153 2999 2167 3013
rect 2233 3019 2247 3033
rect 2293 3007 2307 3021
rect 2313 2999 2327 3013
rect 2333 3007 2347 3021
rect 2353 3019 2367 3033
rect 2373 3027 2387 3041
rect 2453 3039 2467 3053
rect 2393 3019 2407 3033
rect 2473 3027 2487 3041
rect 2413 2999 2427 3013
rect 2513 3019 2527 3033
rect 2533 3027 2547 3041
rect 2553 3019 2567 3033
rect 2613 3019 2627 3033
rect 2573 2999 2587 3013
rect 2813 3076 2827 3090
rect 2653 3019 2667 3033
rect 2693 3007 2707 3021
rect 2713 2999 2727 3013
rect 2733 3007 2747 3021
rect 2953 3076 2967 3090
rect 2853 3019 2867 3033
rect 2893 3019 2907 3033
rect 2973 3047 2987 3061
rect 2953 2982 2967 2996
rect 3053 3039 3067 3053
rect 3033 3019 3047 3033
rect 3073 3019 3087 3033
rect 3113 3019 3127 3033
rect 3133 3027 3147 3041
rect 3153 3039 3167 3053
rect 3173 3027 3187 3041
rect 3213 3039 3227 3053
rect 3193 3019 3207 3033
rect 2813 2950 2827 2964
rect 2953 2944 2967 2958
rect 3313 3076 3327 3090
rect 3233 3019 3247 3033
rect 3453 3076 3467 3090
rect 3353 3019 3367 3033
rect 3393 3019 3407 3033
rect 3473 3047 3487 3061
rect 3453 2982 3467 2996
rect 3313 2950 3327 2964
rect 3453 2944 3467 2958
rect 3553 3076 3567 3090
rect 3693 3076 3707 3090
rect 3593 3019 3607 3033
rect 3633 3019 3647 3033
rect 3713 3047 3727 3061
rect 3693 2982 3707 2996
rect 3773 3039 3787 3053
rect 3753 3019 3767 3033
rect 3793 3019 3807 3033
rect 3873 3019 3887 3033
rect 3893 3027 3907 3041
rect 3913 3019 3927 3033
rect 3973 3019 3987 3033
rect 3993 3027 4007 3041
rect 4013 3019 4027 3033
rect 4033 3019 4047 3033
rect 4053 3027 4067 3041
rect 4073 3019 4087 3033
rect 4133 3019 4147 3033
rect 4153 3027 4167 3041
rect 4233 3039 4247 3053
rect 4273 3073 4287 3087
rect 4173 3019 4187 3033
rect 4253 3027 4267 3041
rect 3853 2999 3867 3013
rect 3953 2999 3967 3013
rect 4093 2999 4107 3013
rect 4193 2999 4207 3013
rect 3553 2950 3567 2964
rect 3693 2944 3707 2958
rect 4433 3076 4447 3090
rect 4573 3076 4587 3090
rect 4413 3047 4427 3061
rect 4273 2993 4287 3007
rect 4293 2999 4307 3013
rect 4333 2999 4347 3013
rect 4353 3007 4367 3021
rect 4313 2979 4327 2993
rect 4433 2982 4447 2996
rect 4493 3019 4507 3033
rect 4533 3019 4547 3033
rect 4733 3073 4747 3087
rect 4633 3019 4647 3033
rect 4653 3027 4667 3041
rect 4673 3019 4687 3033
rect 4693 2999 4707 3013
rect 4733 2993 4747 3007
rect 4433 2944 4447 2958
rect 4573 2950 4587 2964
rect 93 2767 107 2781
rect 33 2739 47 2753
rect 113 2747 127 2761
rect 53 2727 67 2741
rect 133 2739 147 2753
rect 153 2747 167 2761
rect 173 2747 187 2761
rect 193 2739 207 2753
rect 213 2747 227 2761
rect 233 2739 247 2753
rect 253 2747 267 2761
rect 293 2759 307 2773
rect 313 2767 327 2781
rect 333 2759 347 2773
rect 373 2747 387 2761
rect 413 2759 427 2773
rect 493 2767 507 2781
rect 433 2747 447 2761
rect 513 2747 527 2761
rect 533 2739 547 2753
rect 553 2747 567 2761
rect 573 2759 587 2773
rect 593 2767 607 2781
rect 613 2759 627 2773
rect 673 2747 687 2761
rect 693 2739 707 2753
rect 733 2747 747 2761
rect 773 2759 787 2773
rect 793 2767 807 2781
rect 753 2739 767 2753
rect 813 2759 827 2773
rect 853 2747 867 2761
rect 893 2759 907 2773
rect 973 2767 987 2781
rect 1273 2822 1287 2836
rect 1413 2816 1427 2830
rect 913 2747 927 2761
rect 993 2747 1007 2761
rect 1013 2739 1027 2753
rect 1033 2747 1047 2761
rect 1053 2759 1067 2773
rect 1073 2767 1087 2781
rect 1093 2759 1107 2773
rect 1153 2767 1167 2781
rect 1173 2747 1187 2761
rect 1193 2739 1207 2753
rect 1213 2747 1227 2761
rect 1273 2784 1287 2798
rect 1253 2719 1267 2733
rect 1333 2747 1347 2761
rect 1373 2747 1387 2761
rect 1273 2690 1287 2704
rect 1593 2816 1607 2830
rect 1733 2822 1747 2836
rect 1493 2747 1507 2761
rect 1533 2747 1547 2761
rect 1413 2690 1427 2704
rect 1633 2747 1647 2761
rect 1673 2747 1687 2761
rect 1733 2784 1747 2798
rect 1853 2767 1867 2781
rect 1793 2747 1807 2761
rect 1813 2739 1827 2753
rect 1833 2747 1847 2761
rect 1933 2773 1947 2787
rect 1753 2719 1767 2733
rect 1893 2727 1907 2741
rect 1913 2739 1927 2753
rect 1593 2690 1607 2704
rect 1733 2690 1747 2704
rect 1953 2747 1967 2761
rect 1973 2739 1987 2753
rect 1993 2747 2007 2761
rect 1933 2713 1947 2727
rect 2013 2739 2027 2753
rect 2033 2747 2047 2761
rect 2093 2747 2107 2761
rect 2133 2747 2147 2761
rect 2173 2747 2187 2761
rect 2213 2747 2227 2761
rect 2253 2747 2267 2761
rect 2293 2747 2307 2761
rect 2113 2727 2127 2741
rect 2193 2727 2207 2741
rect 2273 2727 2287 2741
rect 2313 2727 2327 2741
rect 2333 2739 2347 2753
rect 2393 2747 2407 2761
rect 2433 2747 2447 2761
rect 2413 2727 2427 2741
rect 2453 2727 2467 2741
rect 2473 2739 2487 2753
rect 2513 2747 2527 2761
rect 2553 2759 2567 2773
rect 2673 2767 2687 2781
rect 2933 2816 2947 2830
rect 3073 2822 3087 2836
rect 2773 2767 2787 2781
rect 2573 2747 2587 2761
rect 2613 2747 2627 2761
rect 2633 2739 2647 2753
rect 2653 2747 2667 2761
rect 2713 2747 2727 2761
rect 2733 2739 2747 2753
rect 2753 2747 2767 2761
rect 2813 2759 2827 2773
rect 2833 2767 2847 2781
rect 2853 2759 2867 2773
rect 2973 2747 2987 2761
rect 3013 2747 3027 2761
rect 3073 2784 3087 2798
rect 3093 2719 3107 2733
rect 2933 2690 2947 2704
rect 3073 2690 3087 2704
rect 3173 2816 3187 2830
rect 3313 2822 3327 2836
rect 3213 2747 3227 2761
rect 3253 2747 3267 2761
rect 3313 2784 3327 2798
rect 3613 2816 3627 2830
rect 3753 2822 3767 2836
rect 3393 2739 3407 2753
rect 3453 2747 3467 2761
rect 3493 2747 3507 2761
rect 3533 2747 3547 2761
rect 3333 2719 3347 2733
rect 3173 2690 3187 2704
rect 3313 2690 3327 2704
rect 3413 2727 3427 2741
rect 3473 2727 3487 2741
rect 3553 2739 3567 2753
rect 3653 2747 3667 2761
rect 3693 2747 3707 2761
rect 3753 2784 3767 2798
rect 3833 2747 3847 2761
rect 3853 2739 3867 2753
rect 3873 2747 3887 2761
rect 3773 2719 3787 2733
rect 3613 2690 3627 2704
rect 3893 2739 3907 2753
rect 3913 2747 3927 2761
rect 3953 2747 3967 2761
rect 4073 2767 4087 2781
rect 4133 2767 4147 2781
rect 4333 2816 4347 2830
rect 4473 2822 4487 2836
rect 3993 2747 4007 2761
rect 4013 2747 4027 2761
rect 3973 2727 3987 2741
rect 4033 2739 4047 2753
rect 4053 2747 4067 2761
rect 3753 2690 3767 2704
rect 4153 2747 4167 2761
rect 4173 2739 4187 2753
rect 4193 2747 4207 2761
rect 4213 2747 4227 2761
rect 4253 2747 4267 2761
rect 4233 2727 4247 2741
rect 4373 2747 4387 2761
rect 4413 2747 4427 2761
rect 4473 2784 4487 2798
rect 4593 2767 4607 2781
rect 4533 2747 4547 2761
rect 4553 2739 4567 2753
rect 4573 2747 4587 2761
rect 4633 2759 4647 2773
rect 4653 2767 4667 2781
rect 4493 2719 4507 2733
rect 4333 2690 4347 2704
rect 4473 2690 4487 2704
rect 4673 2759 4687 2773
rect 113 2547 127 2561
rect 133 2559 147 2573
rect 153 2547 167 2561
rect 13 2519 27 2533
rect 53 2519 67 2533
rect 73 2527 87 2541
rect 173 2539 187 2553
rect 233 2547 247 2561
rect 253 2559 267 2573
rect 33 2499 47 2513
rect 293 2539 307 2553
rect 313 2527 327 2541
rect 353 2539 367 2553
rect 393 2539 407 2553
rect 413 2547 427 2561
rect 433 2559 447 2573
rect 453 2547 467 2561
rect 453 2513 467 2527
rect 493 2593 507 2607
rect 533 2553 547 2567
rect 593 2553 607 2567
rect 493 2527 507 2541
rect 613 2539 627 2553
rect 633 2547 647 2561
rect 653 2539 667 2553
rect 693 2539 707 2553
rect 713 2547 727 2561
rect 513 2519 527 2533
rect 553 2519 567 2533
rect 593 2519 607 2533
rect 533 2499 547 2513
rect 753 2527 767 2541
rect 793 2573 807 2587
rect 773 2519 787 2533
rect 793 2527 807 2541
rect 793 2493 807 2507
rect 833 2527 847 2541
rect 953 2539 967 2553
rect 973 2547 987 2561
rect 993 2539 1007 2553
rect 853 2519 867 2533
rect 893 2519 907 2533
rect 933 2519 947 2533
rect 873 2499 887 2513
rect 1013 2527 1027 2541
rect 1613 2596 1627 2610
rect 1213 2547 1227 2561
rect 1233 2559 1247 2573
rect 1033 2519 1047 2533
rect 1053 2527 1067 2541
rect 1113 2527 1127 2541
rect 1133 2519 1147 2533
rect 1173 2519 1187 2533
rect 1153 2499 1167 2513
rect 1293 2539 1307 2553
rect 1313 2547 1327 2561
rect 1333 2539 1347 2553
rect 1273 2519 1287 2533
rect 1353 2527 1367 2541
rect 1433 2547 1447 2561
rect 1373 2519 1387 2533
rect 1393 2527 1407 2541
rect 1453 2539 1467 2553
rect 1513 2527 1527 2541
rect 1533 2519 1547 2533
rect 1553 2527 1567 2541
rect 1753 2596 1767 2610
rect 1653 2539 1667 2553
rect 1693 2539 1707 2553
rect 1773 2567 1787 2581
rect 1753 2502 1767 2516
rect 1813 2527 1827 2541
rect 1833 2519 1847 2533
rect 1853 2527 1867 2541
rect 1893 2527 1907 2541
rect 2093 2559 2107 2573
rect 1913 2519 1927 2533
rect 1933 2527 1947 2541
rect 1973 2519 1987 2533
rect 2013 2519 2027 2533
rect 2033 2527 2047 2541
rect 2073 2539 2087 2553
rect 1613 2470 1627 2484
rect 1753 2464 1767 2478
rect 1993 2499 2007 2513
rect 2113 2539 2127 2553
rect 2173 2547 2187 2561
rect 2193 2559 2207 2573
rect 2253 2559 2267 2573
rect 2233 2539 2247 2553
rect 2273 2539 2287 2553
rect 2313 2547 2327 2561
rect 2333 2559 2347 2573
rect 2393 2539 2407 2553
rect 2413 2547 2427 2561
rect 2473 2559 2487 2573
rect 2433 2539 2447 2553
rect 2453 2539 2467 2553
rect 2373 2519 2387 2533
rect 2493 2539 2507 2553
rect 2533 2539 2547 2553
rect 2573 2527 2587 2541
rect 2593 2539 2607 2553
rect 2633 2539 2647 2553
rect 2653 2547 2667 2561
rect 2673 2539 2687 2553
rect 2693 2519 2707 2533
rect 2753 2527 2767 2541
rect 2813 2559 2827 2573
rect 2773 2519 2787 2533
rect 2793 2527 2807 2541
rect 2833 2539 2847 2553
rect 2873 2547 2887 2561
rect 2913 2527 2927 2541
rect 2933 2519 2947 2533
rect 2953 2527 2967 2541
rect 2993 2539 3007 2553
rect 3033 2539 3047 2553
rect 3073 2539 3087 2553
rect 3093 2547 3107 2561
rect 3113 2539 3127 2553
rect 3193 2539 3207 2553
rect 3133 2519 3147 2533
rect 3233 2539 3247 2553
rect 3273 2527 3287 2541
rect 3293 2519 3307 2533
rect 3313 2527 3327 2541
rect 3333 2539 3347 2553
rect 3353 2547 3367 2561
rect 3373 2539 3387 2553
rect 3393 2547 3407 2561
rect 3413 2539 3427 2553
rect 3453 2539 3467 2553
rect 3493 2539 3507 2553
rect 3653 2596 3667 2610
rect 3553 2539 3567 2553
rect 3593 2539 3607 2553
rect 3793 2596 3807 2610
rect 3693 2539 3707 2553
rect 3733 2539 3747 2553
rect 3813 2567 3827 2581
rect 3793 2502 3807 2516
rect 4273 2596 4287 2610
rect 3873 2539 3887 2553
rect 3893 2547 3907 2561
rect 3913 2559 3927 2573
rect 3933 2547 3947 2561
rect 3973 2559 3987 2573
rect 3953 2539 3967 2553
rect 3993 2539 4007 2553
rect 4053 2547 4067 2561
rect 4193 2547 4207 2561
rect 4413 2596 4427 2610
rect 4313 2539 4327 2553
rect 4353 2539 4367 2553
rect 3653 2470 3667 2484
rect 3793 2464 3807 2478
rect 4433 2567 4447 2581
rect 4413 2502 4427 2516
rect 4473 2539 4487 2553
rect 4493 2547 4507 2561
rect 4513 2539 4527 2553
rect 4533 2519 4547 2533
rect 4573 2527 4587 2541
rect 4593 2519 4607 2533
rect 4613 2527 4627 2541
rect 4653 2527 4667 2541
rect 4673 2519 4687 2533
rect 4693 2527 4707 2541
rect 4273 2470 4287 2484
rect 4413 2464 4427 2478
rect 73 2307 87 2321
rect 33 2279 47 2293
rect 53 2287 67 2301
rect 93 2287 107 2301
rect 93 2253 107 2267
rect 133 2333 147 2347
rect 133 2287 147 2301
rect 333 2307 347 2321
rect 273 2287 287 2301
rect 313 2287 327 2301
rect 353 2287 367 2301
rect 153 2267 167 2281
rect 173 2259 187 2273
rect 193 2267 207 2281
rect 213 2267 227 2281
rect 233 2259 247 2273
rect 253 2267 267 2281
rect 373 2279 387 2293
rect 573 2287 587 2301
rect 413 2259 427 2273
rect 433 2247 447 2261
rect 453 2259 467 2273
rect 473 2267 487 2281
rect 513 2267 527 2281
rect 533 2259 547 2273
rect 553 2267 567 2281
rect 633 2267 647 2281
rect 653 2259 667 2273
rect 673 2247 687 2261
rect 693 2259 707 2273
rect 713 2247 727 2261
rect 733 2259 747 2273
rect 793 2267 807 2281
rect 813 2279 827 2293
rect 853 2267 867 2281
rect 873 2279 887 2293
rect 893 2287 907 2301
rect 913 2279 927 2293
rect 953 2267 967 2281
rect 1293 2336 1307 2350
rect 1433 2342 1447 2356
rect 993 2279 1007 2293
rect 1073 2287 1087 2301
rect 1173 2287 1187 2301
rect 1013 2267 1027 2281
rect 1093 2267 1107 2281
rect 1113 2259 1127 2273
rect 1133 2267 1147 2281
rect 1193 2267 1207 2281
rect 1213 2259 1227 2273
rect 1233 2267 1247 2281
rect 1333 2267 1347 2281
rect 1373 2267 1387 2281
rect 1433 2304 1447 2318
rect 1633 2336 1647 2350
rect 1773 2342 1787 2356
rect 1513 2287 1527 2301
rect 1453 2239 1467 2253
rect 1533 2267 1547 2281
rect 1553 2259 1567 2273
rect 1573 2267 1587 2281
rect 1293 2210 1307 2224
rect 1433 2210 1447 2224
rect 1673 2267 1687 2281
rect 1713 2267 1727 2281
rect 1773 2304 1787 2318
rect 2093 2336 2107 2350
rect 2233 2342 2247 2356
rect 2013 2287 2027 2301
rect 1853 2259 1867 2273
rect 1793 2239 1807 2253
rect 1633 2210 1647 2224
rect 1773 2210 1787 2224
rect 1873 2247 1887 2261
rect 1913 2259 1927 2273
rect 1953 2267 1967 2281
rect 1933 2247 1947 2261
rect 1973 2259 1987 2273
rect 1993 2267 2007 2281
rect 2133 2267 2147 2281
rect 2173 2267 2187 2281
rect 2233 2304 2247 2318
rect 2513 2307 2527 2321
rect 2493 2287 2507 2301
rect 2533 2287 2547 2301
rect 2313 2267 2327 2281
rect 2253 2239 2267 2253
rect 2093 2210 2107 2224
rect 2233 2210 2247 2224
rect 2333 2259 2347 2273
rect 2353 2247 2367 2261
rect 2373 2259 2387 2273
rect 2413 2267 2427 2281
rect 2553 2279 2567 2293
rect 2433 2259 2447 2273
rect 2453 2247 2467 2261
rect 2473 2259 2487 2273
rect 2593 2267 2607 2281
rect 2733 2342 2747 2356
rect 2873 2336 2887 2350
rect 2633 2279 2647 2293
rect 2653 2267 2667 2281
rect 2733 2304 2747 2318
rect 2713 2239 2727 2253
rect 3273 2342 3287 2356
rect 3413 2336 3427 2350
rect 2793 2267 2807 2281
rect 2833 2267 2847 2281
rect 2733 2210 2747 2224
rect 2953 2287 2967 2301
rect 3053 2287 3067 2301
rect 3193 2287 3207 2301
rect 2973 2267 2987 2281
rect 2993 2259 3007 2273
rect 3013 2267 3027 2281
rect 3073 2267 3087 2281
rect 3093 2259 3107 2273
rect 3113 2267 3127 2281
rect 3133 2267 3147 2281
rect 3153 2259 3167 2273
rect 3173 2267 3187 2281
rect 3273 2304 3287 2318
rect 2873 2210 2887 2224
rect 3253 2239 3267 2253
rect 3333 2267 3347 2281
rect 3373 2267 3387 2281
rect 3273 2210 3287 2224
rect 3493 2287 3507 2301
rect 3513 2267 3527 2281
rect 3533 2259 3547 2273
rect 3553 2267 3567 2281
rect 3593 2267 3607 2281
rect 3633 2267 3647 2281
rect 3673 2267 3687 2281
rect 3613 2247 3627 2261
rect 3653 2247 3667 2261
rect 3413 2210 3427 2224
rect 3773 2313 3787 2327
rect 4113 2336 4127 2350
rect 4253 2342 4267 2356
rect 3733 2273 3747 2287
rect 3773 2279 3787 2293
rect 3793 2287 3807 2301
rect 3713 2259 3727 2273
rect 3813 2279 3827 2293
rect 3953 2293 3967 2307
rect 3853 2267 3867 2281
rect 3873 2259 3887 2273
rect 3893 2267 3907 2281
rect 3913 2259 3927 2273
rect 3933 2267 3947 2281
rect 3933 2233 3947 2247
rect 3973 2267 3987 2281
rect 3993 2259 4007 2273
rect 4013 2267 4027 2281
rect 4033 2259 4047 2273
rect 4053 2267 4067 2281
rect 4153 2267 4167 2281
rect 4193 2267 4207 2281
rect 4253 2304 4267 2318
rect 4273 2239 4287 2253
rect 4113 2210 4127 2224
rect 4253 2210 4267 2224
rect 4353 2342 4367 2356
rect 4493 2336 4507 2350
rect 4353 2304 4367 2318
rect 4333 2239 4347 2253
rect 4413 2267 4427 2281
rect 4453 2267 4467 2281
rect 4353 2210 4367 2224
rect 4613 2287 4627 2301
rect 4553 2267 4567 2281
rect 4573 2259 4587 2273
rect 4593 2267 4607 2281
rect 4653 2279 4667 2293
rect 4673 2287 4687 2301
rect 4493 2210 4507 2224
rect 4693 2279 4707 2293
rect 33 2059 47 2073
rect 73 2059 87 2073
rect 113 2073 127 2087
rect 133 2059 147 2073
rect 153 2067 167 2081
rect 173 2059 187 2073
rect 293 2067 307 2081
rect 313 2079 327 2093
rect 333 2067 347 2081
rect 113 2039 127 2053
rect 213 2047 227 2061
rect 353 2059 367 2073
rect 393 2067 407 2081
rect 413 2079 427 2093
rect 433 2067 447 2081
rect 453 2059 467 2073
rect 693 2067 707 2081
rect 713 2079 727 2093
rect 733 2067 747 2081
rect 113 1993 127 2007
rect 233 2039 247 2053
rect 273 2039 287 2053
rect 253 2019 267 2033
rect 493 2039 507 2053
rect 533 2039 547 2053
rect 553 2047 567 2061
rect 513 2019 527 2033
rect 593 2039 607 2053
rect 633 2039 647 2053
rect 653 2047 667 2061
rect 753 2059 767 2073
rect 833 2059 847 2073
rect 853 2067 867 2081
rect 873 2059 887 2073
rect 1073 2073 1087 2087
rect 1113 2073 1127 2087
rect 1193 2067 1207 2081
rect 1213 2079 1227 2093
rect 1233 2067 1247 2081
rect 613 2019 627 2033
rect 813 2039 827 2053
rect 893 2039 907 2053
rect 933 2039 947 2053
rect 953 2047 967 2061
rect 913 2019 927 2033
rect 993 2039 1007 2053
rect 1033 2039 1047 2053
rect 1053 2047 1067 2061
rect 1013 2019 1027 2033
rect 1093 2039 1107 2053
rect 1133 2039 1147 2053
rect 1153 2047 1167 2061
rect 1253 2059 1267 2073
rect 1113 2019 1127 2033
rect 1293 2093 1307 2107
rect 1313 2079 1327 2093
rect 1293 2059 1307 2073
rect 1273 2033 1287 2047
rect 1333 2059 1347 2073
rect 1373 2053 1387 2067
rect 1353 2013 1367 2027
rect 1393 2047 1407 2061
rect 1433 2093 1447 2107
rect 1413 2039 1427 2053
rect 1433 2047 1447 2061
rect 1473 2047 1487 2061
rect 1493 2039 1507 2053
rect 1513 2047 1527 2061
rect 1533 2047 1547 2061
rect 1553 2039 1567 2053
rect 1573 2047 1587 2061
rect 1653 2059 1667 2073
rect 1673 2067 1687 2081
rect 1693 2059 1707 2073
rect 1713 2067 1727 2081
rect 1733 2079 1747 2093
rect 1753 2067 1767 2081
rect 1833 2079 1847 2093
rect 1773 2059 1787 2073
rect 1813 2059 1827 2073
rect 1633 2039 1647 2053
rect 1473 2013 1487 2027
rect 1853 2059 1867 2073
rect 1933 2059 1947 2073
rect 1953 2067 1967 2081
rect 1973 2059 1987 2073
rect 1993 2059 2007 2073
rect 2013 2067 2027 2081
rect 2033 2059 2047 2073
rect 2133 2059 2147 2073
rect 2153 2067 2167 2081
rect 2173 2059 2187 2073
rect 2213 2067 2227 2081
rect 1913 2039 1927 2053
rect 2053 2039 2067 2053
rect 2113 2039 2127 2053
rect 2353 2067 2367 2081
rect 2393 2047 2407 2061
rect 2413 2039 2427 2053
rect 2433 2047 2447 2061
rect 2493 2059 2507 2073
rect 2513 2047 2527 2061
rect 2573 2079 2587 2093
rect 2553 2059 2567 2073
rect 2593 2059 2607 2073
rect 2633 2067 2647 2081
rect 2693 2047 2707 2061
rect 2873 2116 2887 2130
rect 2713 2039 2727 2053
rect 2733 2047 2747 2061
rect 2753 2047 2767 2061
rect 2773 2039 2787 2053
rect 2793 2047 2807 2061
rect 3013 2116 3027 2130
rect 2913 2059 2927 2073
rect 2953 2059 2967 2073
rect 3033 2087 3047 2101
rect 3013 2022 3027 2036
rect 3413 2116 3427 2130
rect 3093 2059 3107 2073
rect 3113 2067 3127 2081
rect 3133 2079 3147 2093
rect 3153 2067 3167 2081
rect 3193 2079 3207 2093
rect 3173 2059 3187 2073
rect 3213 2059 3227 2073
rect 3273 2059 3287 2073
rect 3293 2067 3307 2081
rect 3313 2059 3327 2073
rect 3333 2067 3347 2081
rect 3353 2059 3367 2073
rect 3553 2116 3567 2130
rect 3753 2116 3767 2130
rect 3453 2059 3467 2073
rect 3493 2059 3507 2073
rect 2873 1990 2887 2004
rect 3013 1984 3027 1998
rect 3573 2087 3587 2101
rect 3553 2022 3567 2036
rect 3613 2059 3627 2073
rect 3633 2067 3647 2081
rect 3653 2059 3667 2073
rect 3673 2039 3687 2053
rect 3893 2116 3907 2130
rect 3793 2059 3807 2073
rect 3833 2059 3847 2073
rect 3413 1990 3427 2004
rect 3553 1984 3567 1998
rect 3913 2087 3927 2101
rect 3893 2022 3907 2036
rect 3753 1990 3767 2004
rect 3893 1984 3907 1998
rect 3993 2116 4007 2130
rect 4133 2116 4147 2130
rect 3973 2087 3987 2101
rect 3993 2022 4007 2036
rect 4053 2059 4067 2073
rect 4093 2059 4107 2073
rect 4213 2059 4227 2073
rect 4233 2067 4247 2081
rect 4253 2059 4267 2073
rect 4273 2067 4287 2081
rect 4313 2079 4327 2093
rect 4573 2116 4587 2130
rect 4713 2116 4727 2130
rect 4293 2059 4307 2073
rect 4333 2067 4347 2081
rect 4413 2079 4427 2093
rect 4493 2079 4507 2093
rect 4553 2087 4567 2101
rect 3993 1984 4007 1998
rect 4133 1990 4147 2004
rect 4393 2059 4407 2073
rect 4433 2059 4447 2073
rect 4473 2059 4487 2073
rect 4513 2059 4527 2073
rect 4573 2022 4587 2036
rect 4633 2059 4647 2073
rect 4673 2059 4687 2073
rect 4573 1984 4587 1998
rect 4713 1990 4727 2004
rect 213 1833 227 1847
rect 193 1807 207 1821
rect 33 1787 47 1801
rect 53 1779 67 1793
rect 73 1787 87 1801
rect 93 1779 107 1793
rect 113 1787 127 1801
rect 133 1787 147 1801
rect 153 1779 167 1793
rect 173 1787 187 1801
rect 193 1773 207 1787
rect 233 1799 247 1813
rect 253 1807 267 1821
rect 373 1827 387 1841
rect 273 1799 287 1813
rect 333 1799 347 1813
rect 353 1807 367 1821
rect 393 1807 407 1821
rect 413 1787 427 1801
rect 433 1779 447 1793
rect 453 1787 467 1801
rect 473 1779 487 1793
rect 493 1787 507 1801
rect 533 1787 547 1801
rect 573 1799 587 1813
rect 593 1787 607 1801
rect 653 1787 667 1801
rect 673 1779 687 1793
rect 693 1787 707 1801
rect 793 1807 807 1821
rect 993 1827 1007 1841
rect 933 1807 947 1821
rect 973 1807 987 1821
rect 1013 1807 1027 1821
rect 733 1787 747 1801
rect 813 1787 827 1801
rect 833 1779 847 1793
rect 853 1787 867 1801
rect 873 1787 887 1801
rect 893 1779 907 1793
rect 913 1787 927 1801
rect 1033 1799 1047 1813
rect 1073 1767 1087 1781
rect 1093 1779 1107 1793
rect 1133 1853 1147 1867
rect 1153 1827 1167 1841
rect 1133 1807 1147 1821
rect 1173 1807 1187 1821
rect 1253 1827 1267 1841
rect 1193 1799 1207 1813
rect 1233 1807 1247 1821
rect 1273 1807 1287 1821
rect 1293 1799 1307 1813
rect 1153 1773 1167 1787
rect 1533 1827 1547 1841
rect 1513 1807 1527 1821
rect 1553 1807 1567 1821
rect 1353 1779 1367 1793
rect 1413 1787 1427 1801
rect 1373 1767 1387 1781
rect 1433 1779 1447 1793
rect 1453 1787 1467 1801
rect 1473 1779 1487 1793
rect 1493 1787 1507 1801
rect 1573 1799 1587 1813
rect 1793 1827 1807 1841
rect 1613 1767 1627 1781
rect 1633 1779 1647 1793
rect 1693 1787 1707 1801
rect 1753 1799 1767 1813
rect 1773 1807 1787 1821
rect 1813 1807 1827 1821
rect 1713 1779 1727 1793
rect 1833 1787 1847 1801
rect 1973 1856 1987 1870
rect 2113 1862 2127 1876
rect 1873 1799 1887 1813
rect 1893 1787 1907 1801
rect 2013 1787 2027 1801
rect 2053 1787 2067 1801
rect 2113 1824 2127 1838
rect 2193 1787 2207 1801
rect 2133 1759 2147 1773
rect 1973 1730 1987 1744
rect 2113 1730 2127 1744
rect 2233 1787 2247 1801
rect 2373 1807 2387 1821
rect 2213 1767 2227 1781
rect 2253 1767 2267 1781
rect 2273 1779 2287 1793
rect 2313 1787 2327 1801
rect 2333 1779 2347 1793
rect 2353 1787 2367 1801
rect 2413 1787 2427 1801
rect 2453 1787 2467 1801
rect 2493 1787 2507 1801
rect 2633 1807 2647 1821
rect 2533 1787 2547 1801
rect 2573 1787 2587 1801
rect 2433 1767 2447 1781
rect 2513 1767 2527 1781
rect 2593 1779 2607 1793
rect 2613 1787 2627 1801
rect 2693 1799 2707 1813
rect 2713 1807 2727 1821
rect 2733 1799 2747 1813
rect 2773 1787 2787 1801
rect 2893 1807 2907 1821
rect 2813 1787 2827 1801
rect 2833 1787 2847 1801
rect 2793 1767 2807 1781
rect 2853 1779 2867 1793
rect 2873 1787 2887 1801
rect 3113 1862 3127 1876
rect 3253 1856 3267 1870
rect 2933 1767 2947 1781
rect 2953 1779 2967 1793
rect 3013 1787 3027 1801
rect 3053 1787 3067 1801
rect 3033 1767 3047 1781
rect 3113 1824 3127 1838
rect 3093 1759 3107 1773
rect 3173 1787 3187 1801
rect 3213 1787 3227 1801
rect 3113 1730 3127 1744
rect 3533 1862 3547 1876
rect 3673 1856 3687 1870
rect 3373 1807 3387 1821
rect 3313 1787 3327 1801
rect 3333 1779 3347 1793
rect 3353 1787 3367 1801
rect 3413 1799 3427 1813
rect 3433 1807 3447 1821
rect 3253 1730 3267 1744
rect 3453 1799 3467 1813
rect 3533 1824 3547 1838
rect 3513 1759 3527 1773
rect 3593 1787 3607 1801
rect 3633 1787 3647 1801
rect 3533 1730 3547 1744
rect 3733 1787 3747 1801
rect 3773 1787 3787 1801
rect 3833 1799 3847 1813
rect 3853 1807 3867 1821
rect 3673 1730 3687 1744
rect 3873 1799 3887 1813
rect 3913 1853 3927 1867
rect 3913 1807 3927 1821
rect 4013 1807 4027 1821
rect 3933 1787 3947 1801
rect 3913 1773 3927 1787
rect 3953 1779 3967 1793
rect 3973 1787 3987 1801
rect 4033 1787 4047 1801
rect 4053 1779 4067 1793
rect 4073 1787 4087 1801
rect 4113 1787 4127 1801
rect 4093 1767 4107 1781
rect 4473 1862 4487 1876
rect 4613 1856 4627 1870
rect 4153 1779 4167 1793
rect 4213 1779 4227 1793
rect 4233 1767 4247 1781
rect 4253 1779 4267 1793
rect 4273 1767 4287 1781
rect 4293 1779 4307 1793
rect 4313 1787 4327 1801
rect 4373 1787 4387 1801
rect 4413 1787 4427 1801
rect 4393 1767 4407 1781
rect 4473 1824 4487 1838
rect 4453 1759 4467 1773
rect 4533 1787 4547 1801
rect 4573 1787 4587 1801
rect 4473 1730 4487 1744
rect 4693 1799 4707 1813
rect 4713 1807 4727 1821
rect 4733 1799 4747 1813
rect 4613 1730 4627 1744
rect 33 1587 47 1601
rect 53 1599 67 1613
rect 93 1579 107 1593
rect 113 1587 127 1601
rect 133 1599 147 1613
rect 153 1587 167 1601
rect 173 1559 187 1573
rect 213 1559 227 1573
rect 233 1567 247 1581
rect 193 1539 207 1553
rect 273 1613 287 1627
rect 273 1567 287 1581
rect 293 1559 307 1573
rect 313 1567 327 1581
rect 393 1579 407 1593
rect 413 1587 427 1601
rect 433 1579 447 1593
rect 473 1579 487 1593
rect 373 1559 387 1573
rect 273 1533 287 1547
rect 513 1579 527 1593
rect 553 1587 567 1601
rect 573 1599 587 1613
rect 693 1587 707 1601
rect 713 1599 727 1613
rect 733 1587 747 1601
rect 593 1559 607 1573
rect 633 1559 647 1573
rect 653 1567 667 1581
rect 753 1579 767 1593
rect 893 1587 907 1601
rect 913 1599 927 1613
rect 933 1587 947 1601
rect 1073 1613 1087 1627
rect 1253 1633 1267 1647
rect 613 1539 627 1553
rect 793 1559 807 1573
rect 833 1559 847 1573
rect 853 1567 867 1581
rect 953 1579 967 1593
rect 813 1539 827 1553
rect 993 1559 1007 1573
rect 1033 1559 1047 1573
rect 1053 1567 1067 1581
rect 1013 1539 1027 1553
rect 1133 1579 1147 1593
rect 1153 1587 1167 1601
rect 1173 1579 1187 1593
rect 1113 1559 1127 1573
rect 1093 1533 1107 1547
rect 1193 1559 1207 1573
rect 1233 1559 1247 1573
rect 1253 1567 1267 1581
rect 1213 1539 1227 1553
rect 1293 1587 1307 1601
rect 1313 1599 1327 1613
rect 1333 1587 1347 1601
rect 1353 1579 1367 1593
rect 1413 1587 1427 1601
rect 1433 1599 1447 1613
rect 1293 1553 1307 1567
rect 1553 1587 1567 1601
rect 1573 1599 1587 1613
rect 1593 1587 1607 1601
rect 1453 1559 1467 1573
rect 1493 1559 1507 1573
rect 1513 1567 1527 1581
rect 1613 1579 1627 1593
rect 1473 1539 1487 1553
rect 1653 1559 1667 1573
rect 1693 1559 1707 1573
rect 1713 1567 1727 1581
rect 1753 1579 1767 1593
rect 1773 1587 1787 1601
rect 1793 1579 1807 1593
rect 1873 1579 1887 1593
rect 1893 1587 1907 1601
rect 1913 1599 1927 1613
rect 1933 1587 1947 1601
rect 1953 1599 1967 1613
rect 1973 1587 1987 1601
rect 1673 1539 1687 1553
rect 1813 1559 1827 1573
rect 2033 1593 2047 1607
rect 2013 1559 2027 1573
rect 2053 1559 2067 1573
rect 2073 1567 2087 1581
rect 1993 1533 2007 1547
rect 2033 1539 2047 1553
rect 2093 1533 2107 1547
rect 2133 1593 2147 1607
rect 2153 1579 2167 1593
rect 2173 1587 2187 1601
rect 2213 1599 2227 1613
rect 2313 1636 2327 1650
rect 2453 1636 2467 1650
rect 2293 1607 2307 1621
rect 2193 1579 2207 1593
rect 2233 1587 2247 1601
rect 2133 1559 2147 1573
rect 2313 1542 2327 1556
rect 2373 1579 2387 1593
rect 2413 1579 2427 1593
rect 2553 1579 2567 1593
rect 2573 1587 2587 1601
rect 2593 1579 2607 1593
rect 2633 1579 2647 1593
rect 2533 1559 2547 1573
rect 2653 1567 2667 1581
rect 2313 1504 2327 1518
rect 2453 1510 2467 1524
rect 2733 1599 2747 1613
rect 2693 1579 2707 1593
rect 2713 1579 2727 1593
rect 2753 1579 2767 1593
rect 2793 1587 2807 1601
rect 2813 1599 2827 1613
rect 2833 1587 2847 1601
rect 2933 1599 2947 1613
rect 2853 1579 2867 1593
rect 2913 1579 2927 1593
rect 2953 1579 2967 1593
rect 2993 1587 3007 1601
rect 3013 1599 3027 1613
rect 3053 1587 3067 1601
rect 3073 1599 3087 1613
rect 3093 1579 3107 1593
rect 3113 1587 3127 1601
rect 3133 1579 3147 1593
rect 3153 1559 3167 1573
rect 3193 1567 3207 1581
rect 3213 1559 3227 1573
rect 3233 1567 3247 1581
rect 3293 1567 3307 1581
rect 3493 1636 3507 1650
rect 3313 1559 3327 1573
rect 3333 1567 3347 1581
rect 3373 1593 3387 1607
rect 3393 1579 3407 1593
rect 3413 1587 3427 1601
rect 3433 1579 3447 1593
rect 3373 1559 3387 1573
rect 3633 1636 3647 1650
rect 3533 1579 3547 1593
rect 3573 1579 3587 1593
rect 3373 1513 3387 1527
rect 3653 1607 3667 1621
rect 3633 1542 3647 1556
rect 3693 1599 3707 1613
rect 3713 1587 3727 1601
rect 3773 1587 3787 1601
rect 3793 1599 3807 1613
rect 3493 1510 3507 1524
rect 3633 1504 3647 1518
rect 3853 1579 3867 1593
rect 3873 1587 3887 1601
rect 3933 1599 3947 1613
rect 4013 1599 4027 1613
rect 4073 1599 4087 1613
rect 3893 1579 3907 1593
rect 3913 1579 3927 1593
rect 3833 1559 3847 1573
rect 3953 1579 3967 1593
rect 3993 1579 4007 1593
rect 4033 1579 4047 1593
rect 4093 1587 4107 1601
rect 4133 1587 4147 1601
rect 4153 1599 4167 1613
rect 4173 1587 4187 1601
rect 4213 1613 4227 1627
rect 4193 1579 4207 1593
rect 4253 1599 4267 1613
rect 4233 1579 4247 1593
rect 4213 1553 4227 1567
rect 4273 1579 4287 1593
rect 4313 1587 4327 1601
rect 4333 1599 4347 1613
rect 4353 1587 4367 1601
rect 4413 1599 4427 1613
rect 4373 1579 4387 1593
rect 4433 1587 4447 1601
rect 4473 1599 4487 1613
rect 4493 1587 4507 1601
rect 4553 1587 4567 1601
rect 4573 1599 4587 1613
rect 4593 1579 4607 1593
rect 4613 1587 4627 1601
rect 4673 1613 4687 1627
rect 4633 1579 4647 1593
rect 4653 1559 4667 1573
rect 4653 1513 4667 1527
rect 4693 1567 4707 1581
rect 4713 1559 4727 1573
rect 4733 1567 4747 1581
rect 133 1347 147 1361
rect 113 1327 127 1341
rect 153 1327 167 1341
rect 193 1353 207 1367
rect 33 1307 47 1321
rect 173 1319 187 1333
rect 53 1299 67 1313
rect 73 1287 87 1301
rect 93 1299 107 1313
rect 233 1347 247 1361
rect 213 1327 227 1341
rect 253 1327 267 1341
rect 293 1353 307 1367
rect 273 1319 287 1333
rect 213 1293 227 1307
rect 333 1319 347 1333
rect 353 1327 367 1341
rect 293 1273 307 1287
rect 373 1319 387 1333
rect 473 1353 487 1367
rect 453 1327 467 1341
rect 393 1307 407 1321
rect 413 1299 427 1313
rect 433 1307 447 1321
rect 653 1327 667 1341
rect 753 1327 767 1341
rect 473 1293 487 1307
rect 493 1299 507 1313
rect 513 1287 527 1301
rect 533 1299 547 1313
rect 553 1307 567 1321
rect 593 1307 607 1321
rect 613 1299 627 1313
rect 633 1307 647 1321
rect 693 1307 707 1321
rect 713 1299 727 1313
rect 733 1307 747 1321
rect 793 1307 807 1321
rect 833 1319 847 1333
rect 853 1307 867 1321
rect 913 1319 927 1333
rect 933 1327 947 1341
rect 953 1319 967 1333
rect 973 1319 987 1333
rect 993 1327 1007 1341
rect 1113 1347 1127 1361
rect 1013 1319 1027 1333
rect 1073 1319 1087 1333
rect 1093 1327 1107 1341
rect 1133 1327 1147 1341
rect 1173 1299 1187 1313
rect 1233 1307 1247 1321
rect 1253 1319 1267 1333
rect 1193 1287 1207 1301
rect 1373 1327 1387 1341
rect 1293 1307 1307 1321
rect 1313 1307 1327 1321
rect 1333 1299 1347 1313
rect 1353 1307 1367 1321
rect 1433 1373 1447 1387
rect 1433 1327 1447 1341
rect 1453 1307 1467 1321
rect 1433 1293 1447 1307
rect 1473 1299 1487 1313
rect 1493 1307 1507 1321
rect 1513 1319 1527 1333
rect 1533 1327 1547 1341
rect 1553 1319 1567 1333
rect 1653 1327 1667 1341
rect 1593 1307 1607 1321
rect 1613 1299 1627 1313
rect 1633 1307 1647 1321
rect 1693 1319 1707 1333
rect 1713 1327 1727 1341
rect 1733 1319 1747 1333
rect 1893 1347 1907 1361
rect 1873 1327 1887 1341
rect 1913 1327 1927 1341
rect 1773 1299 1787 1313
rect 1793 1287 1807 1301
rect 1813 1299 1827 1313
rect 1833 1307 1847 1321
rect 1933 1319 1947 1333
rect 2033 1327 2047 1341
rect 1973 1307 1987 1321
rect 1993 1299 2007 1313
rect 2013 1307 2027 1321
rect 2153 1347 2167 1361
rect 2133 1327 2147 1341
rect 2173 1327 2187 1341
rect 2193 1319 2207 1333
rect 2233 1319 2247 1333
rect 2253 1327 2267 1341
rect 2073 1287 2087 1301
rect 2093 1299 2107 1313
rect 2273 1319 2287 1333
rect 2333 1307 2347 1321
rect 2313 1287 2327 1301
rect 2433 1319 2447 1333
rect 2453 1327 2467 1341
rect 2373 1299 2387 1313
rect 2473 1319 2487 1333
rect 2893 1376 2907 1390
rect 3033 1382 3047 1396
rect 2493 1287 2507 1301
rect 2513 1299 2527 1313
rect 2573 1307 2587 1321
rect 2693 1327 2707 1341
rect 2613 1307 2627 1321
rect 2633 1307 2647 1321
rect 2653 1299 2667 1313
rect 2673 1307 2687 1321
rect 2753 1307 2767 1321
rect 2773 1299 2787 1313
rect 2793 1307 2807 1321
rect 2813 1299 2827 1313
rect 2833 1307 2847 1321
rect 2933 1307 2947 1321
rect 2973 1307 2987 1321
rect 3033 1344 3047 1358
rect 3313 1376 3327 1390
rect 3453 1382 3467 1396
rect 3113 1307 3127 1321
rect 3053 1279 3067 1293
rect 2893 1250 2907 1264
rect 3033 1250 3047 1264
rect 3153 1307 3167 1321
rect 3193 1307 3207 1321
rect 3133 1287 3147 1301
rect 3213 1299 3227 1313
rect 3233 1287 3247 1301
rect 3253 1299 3267 1313
rect 3353 1307 3367 1321
rect 3393 1307 3407 1321
rect 3453 1344 3467 1358
rect 3533 1299 3547 1313
rect 3593 1307 3607 1321
rect 3633 1307 3647 1321
rect 3673 1307 3687 1321
rect 3713 1307 3727 1321
rect 3833 1382 3847 1396
rect 3973 1376 3987 1390
rect 3473 1279 3487 1293
rect 3313 1250 3327 1264
rect 3453 1250 3467 1264
rect 3553 1287 3567 1301
rect 3613 1287 3627 1301
rect 3693 1287 3707 1301
rect 3733 1287 3747 1301
rect 3753 1299 3767 1313
rect 3833 1344 3847 1358
rect 3813 1279 3827 1293
rect 3893 1307 3907 1321
rect 3933 1307 3947 1321
rect 3833 1250 3847 1264
rect 4093 1327 4107 1341
rect 4033 1307 4047 1321
rect 4053 1299 4067 1313
rect 4073 1307 4087 1321
rect 4133 1319 4147 1333
rect 4153 1327 4167 1341
rect 3973 1250 3987 1264
rect 4173 1319 4187 1333
rect 4233 1307 4247 1321
rect 4273 1307 4287 1321
rect 4313 1319 4327 1333
rect 4333 1327 4347 1341
rect 4353 1319 4367 1333
rect 4393 1327 4407 1341
rect 4493 1327 4507 1341
rect 4413 1307 4427 1321
rect 4433 1299 4447 1313
rect 4453 1307 4467 1321
rect 4513 1307 4527 1321
rect 4533 1299 4547 1313
rect 4553 1307 4567 1321
rect 4573 1307 4587 1321
rect 4613 1307 4627 1321
rect 4593 1287 4607 1301
rect 4653 1287 4667 1301
rect 4673 1299 4687 1313
rect 4733 1299 4747 1313
rect 4753 1287 4767 1301
rect 53 1099 67 1113
rect 73 1107 87 1121
rect 93 1099 107 1113
rect 113 1099 127 1113
rect 133 1107 147 1121
rect 293 1133 307 1147
rect 153 1099 167 1113
rect 33 1079 47 1093
rect 173 1079 187 1093
rect 213 1079 227 1093
rect 253 1079 267 1093
rect 273 1087 287 1101
rect 313 1107 327 1121
rect 333 1119 347 1133
rect 353 1107 367 1121
rect 473 1153 487 1167
rect 373 1099 387 1113
rect 233 1059 247 1073
rect 293 1073 307 1087
rect 413 1079 427 1093
rect 453 1079 467 1093
rect 473 1087 487 1101
rect 433 1059 447 1073
rect 513 1107 527 1121
rect 533 1119 547 1133
rect 553 1107 567 1121
rect 573 1099 587 1113
rect 513 1073 527 1087
rect 633 1087 647 1101
rect 653 1079 667 1093
rect 673 1087 687 1101
rect 713 1099 727 1113
rect 733 1087 747 1101
rect 773 1099 787 1113
rect 853 1113 867 1127
rect 813 1087 827 1101
rect 833 1079 847 1093
rect 873 1079 887 1093
rect 853 1059 867 1073
rect 933 1099 947 1113
rect 953 1107 967 1121
rect 973 1099 987 1113
rect 993 1099 1007 1113
rect 1013 1107 1027 1121
rect 1033 1099 1047 1113
rect 1133 1099 1147 1113
rect 1153 1107 1167 1121
rect 1173 1099 1187 1113
rect 913 1079 927 1093
rect 1053 1079 1067 1093
rect 1113 1079 1127 1093
rect 1213 1087 1227 1101
rect 1233 1079 1247 1093
rect 1253 1087 1267 1101
rect 1293 1099 1307 1113
rect 893 1033 907 1047
rect 1313 1087 1327 1101
rect 1353 1099 1367 1113
rect 1373 1087 1387 1101
rect 1393 1079 1407 1093
rect 1413 1087 1427 1101
rect 1473 1099 1487 1113
rect 1493 1107 1507 1121
rect 1533 1087 1547 1101
rect 1573 1133 1587 1147
rect 1553 1079 1567 1093
rect 1573 1087 1587 1101
rect 1613 1087 1627 1101
rect 1633 1079 1647 1093
rect 1653 1087 1667 1101
rect 1673 1079 1687 1093
rect 1713 1079 1727 1093
rect 1733 1087 1747 1101
rect 1793 1087 1807 1101
rect 1613 1033 1627 1047
rect 1693 1059 1707 1073
rect 1813 1079 1827 1093
rect 1833 1087 1847 1101
rect 1853 1079 1867 1093
rect 1893 1079 1907 1093
rect 1913 1087 1927 1101
rect 1953 1087 1967 1101
rect 1873 1059 1887 1073
rect 1973 1079 1987 1093
rect 1993 1087 2007 1101
rect 2053 1099 2067 1113
rect 2073 1107 2087 1121
rect 2093 1099 2107 1113
rect 2113 1107 2127 1121
rect 2133 1099 2147 1113
rect 2213 1113 2227 1127
rect 2173 1087 2187 1101
rect 2193 1079 2207 1093
rect 2233 1079 2247 1093
rect 2213 1059 2227 1073
rect 2273 1087 2287 1101
rect 2333 1107 2347 1121
rect 2353 1119 2367 1133
rect 2373 1107 2387 1121
rect 2293 1079 2307 1093
rect 2313 1087 2327 1101
rect 2393 1099 2407 1113
rect 2453 1107 2467 1121
rect 2473 1119 2487 1133
rect 2273 1053 2287 1067
rect 2513 1087 2527 1101
rect 2813 1156 2827 1170
rect 2533 1079 2547 1093
rect 2553 1087 2567 1101
rect 2593 1099 2607 1113
rect 2613 1107 2627 1121
rect 2633 1099 2647 1113
rect 2653 1107 2667 1121
rect 2673 1099 2687 1113
rect 2693 1099 2707 1113
rect 2733 1099 2747 1113
rect 2953 1156 2967 1170
rect 2853 1099 2867 1113
rect 2893 1099 2907 1113
rect 2973 1127 2987 1141
rect 2953 1062 2967 1076
rect 3013 1087 3027 1101
rect 3033 1079 3047 1093
rect 3053 1087 3067 1101
rect 3133 1099 3147 1113
rect 3153 1107 3167 1121
rect 3173 1099 3187 1113
rect 3213 1099 3227 1113
rect 3253 1099 3267 1113
rect 3333 1099 3347 1113
rect 3113 1079 3127 1093
rect 2813 1030 2827 1044
rect 2953 1024 2967 1038
rect 3373 1099 3387 1113
rect 3393 1099 3407 1113
rect 3433 1099 3447 1113
rect 3493 1107 3507 1121
rect 3633 1107 3647 1121
rect 3693 1107 3707 1121
rect 3833 1107 3847 1121
rect 3873 1099 3887 1113
rect 4073 1156 4087 1170
rect 3913 1099 3927 1113
rect 3953 1087 3967 1101
rect 4213 1156 4227 1170
rect 4053 1127 4067 1141
rect 3973 1079 3987 1093
rect 3993 1087 4007 1101
rect 4073 1062 4087 1076
rect 4133 1099 4147 1113
rect 4173 1099 4187 1113
rect 4273 1087 4287 1101
rect 4293 1079 4307 1093
rect 4313 1087 4327 1101
rect 4353 1099 4367 1113
rect 4373 1107 4387 1121
rect 4393 1099 4407 1113
rect 4073 1024 4087 1038
rect 4213 1030 4227 1044
rect 4413 1079 4427 1093
rect 4473 1087 4487 1101
rect 4493 1079 4507 1093
rect 4513 1087 4527 1101
rect 4533 1099 4547 1113
rect 4553 1107 4567 1121
rect 4573 1099 4587 1113
rect 4593 1079 4607 1093
rect 4633 1079 4647 1093
rect 4673 1079 4687 1093
rect 4693 1087 4707 1101
rect 4653 1059 4667 1073
rect 33 839 47 853
rect 53 847 67 861
rect 73 839 87 853
rect 113 827 127 841
rect 133 839 147 853
rect 213 847 227 861
rect 173 827 187 841
rect 233 827 247 841
rect 253 819 267 833
rect 273 827 287 841
rect 313 827 327 841
rect 333 819 347 833
rect 353 827 367 841
rect 373 819 387 833
rect 393 827 407 841
rect 433 827 447 841
rect 473 827 487 841
rect 733 867 747 881
rect 713 847 727 861
rect 753 847 767 861
rect 493 807 507 821
rect 513 819 527 833
rect 573 819 587 833
rect 633 827 647 841
rect 773 839 787 853
rect 593 807 607 821
rect 653 819 667 833
rect 673 807 687 821
rect 693 819 707 833
rect 833 827 847 841
rect 853 839 867 853
rect 893 827 907 841
rect 913 839 927 853
rect 933 847 947 861
rect 1053 867 1067 881
rect 953 839 967 853
rect 1013 839 1027 853
rect 1033 847 1047 861
rect 1073 847 1087 861
rect 1153 847 1167 861
rect 1253 867 1267 881
rect 1093 827 1107 841
rect 1113 819 1127 833
rect 1133 827 1147 841
rect 1213 839 1227 853
rect 1233 847 1247 861
rect 1273 847 1287 861
rect 1613 933 1627 947
rect 1573 873 1587 887
rect 1413 847 1427 861
rect 1293 807 1307 821
rect 1313 819 1327 833
rect 1353 827 1367 841
rect 1373 819 1387 833
rect 1393 827 1407 841
rect 1473 839 1487 853
rect 1493 847 1507 861
rect 1513 839 1527 853
rect 1533 839 1547 853
rect 1553 847 1567 861
rect 1593 853 1607 867
rect 1573 839 1587 853
rect 1633 847 1647 861
rect 1653 827 1667 841
rect 1633 813 1647 827
rect 1673 819 1687 833
rect 1693 827 1707 841
rect 1713 827 1727 841
rect 1753 839 1767 853
rect 1773 827 1787 841
rect 1893 839 1907 853
rect 1913 847 1927 861
rect 1833 819 1847 833
rect 1853 807 1867 821
rect 1933 839 1947 853
rect 2073 867 2087 881
rect 2033 839 2047 853
rect 2053 847 2067 861
rect 2093 847 2107 861
rect 1953 807 1967 821
rect 1973 819 1987 833
rect 2233 847 2247 861
rect 2113 807 2127 821
rect 2133 819 2147 833
rect 2173 827 2187 841
rect 2193 819 2207 833
rect 2213 827 2227 841
rect 2293 827 2307 841
rect 2453 867 2467 881
rect 2433 847 2447 861
rect 2473 847 2487 861
rect 2593 867 2607 881
rect 2493 839 2507 853
rect 2553 839 2567 853
rect 2573 847 2587 861
rect 2613 847 2627 861
rect 2313 819 2327 833
rect 2333 807 2347 821
rect 2353 819 2367 833
rect 2373 807 2387 821
rect 2393 819 2407 833
rect 2633 819 2647 833
rect 2653 807 2667 821
rect 2673 819 2687 833
rect 2693 827 2707 841
rect 2753 839 2767 853
rect 2773 847 2787 861
rect 2793 839 2807 853
rect 2833 827 2847 841
rect 2853 819 2867 833
rect 2873 827 2887 841
rect 2893 819 2907 833
rect 2913 827 2927 841
rect 2953 819 2967 833
rect 3013 827 3027 841
rect 3053 827 3067 841
rect 3093 827 3107 841
rect 3133 827 3147 841
rect 3433 902 3447 916
rect 3573 896 3587 910
rect 3273 847 3287 861
rect 2973 807 2987 821
rect 3033 807 3047 821
rect 3113 807 3127 821
rect 3153 807 3167 821
rect 3173 819 3187 833
rect 3213 827 3227 841
rect 3233 819 3247 833
rect 3253 827 3267 841
rect 3313 839 3327 853
rect 3333 847 3347 861
rect 3353 839 3367 853
rect 3433 864 3447 878
rect 3413 799 3427 813
rect 3493 827 3507 841
rect 3533 827 3547 841
rect 3433 770 3447 784
rect 3753 896 3767 910
rect 3893 902 3907 916
rect 3633 827 3647 841
rect 3673 827 3687 841
rect 3573 770 3587 784
rect 3793 827 3807 841
rect 3833 827 3847 841
rect 3893 864 3907 878
rect 4093 902 4107 916
rect 4233 896 4247 910
rect 3973 847 3987 861
rect 3913 799 3927 813
rect 3993 827 4007 841
rect 4013 819 4027 833
rect 4033 827 4047 841
rect 4093 864 4107 878
rect 3753 770 3767 784
rect 4073 799 4087 813
rect 4153 827 4167 841
rect 4193 827 4207 841
rect 3893 770 3907 784
rect 4093 770 4107 784
rect 4233 770 4247 784
rect 4333 896 4347 910
rect 4473 902 4487 916
rect 4373 827 4387 841
rect 4413 827 4427 841
rect 4473 864 4487 878
rect 4593 847 4607 861
rect 4693 847 4707 861
rect 4533 827 4547 841
rect 4553 819 4567 833
rect 4573 827 4587 841
rect 4633 827 4647 841
rect 4493 799 4507 813
rect 4653 819 4667 833
rect 4673 827 4687 841
rect 4333 770 4347 784
rect 4473 770 4487 784
rect 53 639 67 653
rect 33 619 47 633
rect 73 619 87 633
rect 113 619 127 633
rect 133 627 147 641
rect 153 639 167 653
rect 173 627 187 641
rect 193 639 207 653
rect 213 627 227 641
rect 273 619 287 633
rect 293 627 307 641
rect 313 639 327 653
rect 333 627 347 641
rect 353 599 367 613
rect 393 599 407 613
rect 413 607 427 621
rect 493 619 507 633
rect 513 627 527 641
rect 533 619 547 633
rect 573 619 587 633
rect 373 579 387 593
rect 473 599 487 613
rect 613 619 627 633
rect 673 619 687 633
rect 693 627 707 641
rect 713 619 727 633
rect 753 619 767 633
rect 653 599 667 613
rect 793 619 807 633
rect 813 619 827 633
rect 853 607 867 621
rect 873 619 887 633
rect 913 619 927 633
rect 933 627 947 641
rect 953 619 967 633
rect 1053 619 1067 633
rect 1073 627 1087 641
rect 1093 619 1107 633
rect 1133 619 1147 633
rect 1153 627 1167 641
rect 1173 627 1187 641
rect 1193 639 1207 653
rect 1213 627 1227 641
rect 1233 619 1247 633
rect 1293 627 1307 641
rect 1313 639 1327 653
rect 973 599 987 613
rect 1033 599 1047 613
rect 1333 619 1347 633
rect 1353 627 1367 641
rect 1373 619 1387 633
rect 1433 619 1447 633
rect 1453 627 1467 641
rect 1473 619 1487 633
rect 1553 619 1567 633
rect 1573 627 1587 641
rect 1593 639 1607 653
rect 1613 627 1627 641
rect 1633 627 1647 641
rect 1653 639 1667 653
rect 1673 627 1687 641
rect 1693 619 1707 633
rect 1393 599 1407 613
rect 1493 599 1507 613
rect 1733 599 1747 613
rect 1773 599 1787 613
rect 1793 607 1807 621
rect 1833 619 1847 633
rect 1853 627 1867 641
rect 1893 633 1907 647
rect 1873 619 1887 633
rect 1753 579 1767 593
rect 1893 599 1907 613
rect 1893 553 1907 567
rect 2153 673 2167 687
rect 1953 619 1967 633
rect 1973 627 1987 641
rect 1993 639 2007 653
rect 2013 627 2027 641
rect 2033 619 2047 633
rect 2053 627 2067 641
rect 2073 619 2087 633
rect 2093 599 2107 613
rect 2233 633 2247 647
rect 2153 607 2167 621
rect 2113 573 2127 587
rect 2173 599 2187 613
rect 2213 599 2227 613
rect 2193 579 2207 593
rect 2213 553 2227 567
rect 2273 619 2287 633
rect 2293 627 2307 641
rect 2313 619 2327 633
rect 2333 619 2347 633
rect 2353 627 2367 641
rect 2373 619 2387 633
rect 2833 676 2847 690
rect 2653 627 2667 641
rect 2673 639 2687 653
rect 2253 599 2267 613
rect 2393 599 2407 613
rect 2433 599 2447 613
rect 2473 599 2487 613
rect 2493 607 2507 621
rect 2453 579 2467 593
rect 2533 599 2547 613
rect 2573 599 2587 613
rect 2593 607 2607 621
rect 2553 579 2567 593
rect 2693 599 2707 613
rect 2733 599 2747 613
rect 2753 607 2767 621
rect 2713 579 2727 593
rect 2973 676 2987 690
rect 2873 619 2887 633
rect 2913 619 2927 633
rect 2993 647 3007 661
rect 2973 582 2987 596
rect 3033 619 3047 633
rect 3053 627 3067 641
rect 3133 639 3147 653
rect 3073 619 3087 633
rect 3153 627 3167 641
rect 3193 639 3207 653
rect 3213 627 3227 641
rect 3093 599 3107 613
rect 2833 550 2847 564
rect 2973 544 2987 558
rect 3373 627 3387 641
rect 3393 639 3407 653
rect 3253 599 3267 613
rect 3293 599 3307 613
rect 3313 607 3327 621
rect 3273 579 3287 593
rect 3433 607 3447 621
rect 3633 676 3647 690
rect 3453 599 3467 613
rect 3473 607 3487 621
rect 3533 619 3547 633
rect 3553 627 3567 641
rect 3573 619 3587 633
rect 3513 599 3527 613
rect 3773 676 3787 690
rect 4053 676 4067 690
rect 3673 619 3687 633
rect 3713 619 3727 633
rect 3793 647 3807 661
rect 3773 582 3787 596
rect 3833 619 3847 633
rect 3853 627 3867 641
rect 3873 619 3887 633
rect 3893 599 3907 613
rect 3953 607 3967 621
rect 4193 676 4207 690
rect 4033 647 4047 661
rect 3973 599 3987 613
rect 3993 607 4007 621
rect 3633 550 3647 564
rect 3773 544 3787 558
rect 4053 582 4067 596
rect 4113 619 4127 633
rect 4153 619 4167 633
rect 4553 676 4567 690
rect 4253 607 4267 621
rect 4273 599 4287 613
rect 4293 607 4307 621
rect 4333 607 4347 621
rect 4353 599 4367 613
rect 4373 607 4387 621
rect 4453 619 4467 633
rect 4473 627 4487 641
rect 4493 619 4507 633
rect 4433 599 4447 613
rect 4053 544 4067 558
rect 4193 550 4207 564
rect 4693 676 4707 690
rect 4593 619 4607 633
rect 4633 619 4647 633
rect 4713 647 4727 661
rect 4693 582 4707 596
rect 4553 550 4567 564
rect 4693 544 4707 558
rect 233 393 247 407
rect 13 359 27 373
rect 33 367 47 381
rect 53 359 67 373
rect 93 359 107 373
rect 113 367 127 381
rect 133 359 147 373
rect 193 359 207 373
rect 213 367 227 381
rect 233 359 247 373
rect 273 359 287 373
rect 293 367 307 381
rect 253 333 267 347
rect 313 359 327 373
rect 353 347 367 361
rect 373 359 387 373
rect 413 393 427 407
rect 413 347 427 361
rect 453 359 467 373
rect 473 367 487 381
rect 573 387 587 401
rect 493 359 507 373
rect 533 359 547 373
rect 553 367 567 381
rect 593 367 607 381
rect 633 347 647 361
rect 653 339 667 353
rect 673 347 687 361
rect 433 293 447 307
rect 693 339 707 353
rect 713 347 727 361
rect 753 347 767 361
rect 793 347 807 361
rect 833 359 847 373
rect 853 367 867 381
rect 773 327 787 341
rect 873 359 887 373
rect 893 359 907 373
rect 913 367 927 381
rect 933 359 947 373
rect 993 359 1007 373
rect 1013 367 1027 381
rect 1033 359 1047 373
rect 1073 359 1087 373
rect 1093 367 1107 381
rect 1113 359 1127 373
rect 1313 367 1327 381
rect 1153 347 1167 361
rect 1173 339 1187 353
rect 1193 347 1207 361
rect 1213 339 1227 353
rect 1233 347 1247 361
rect 1253 347 1267 361
rect 1273 339 1287 353
rect 1293 347 1307 361
rect 1373 347 1387 361
rect 1493 367 1507 381
rect 1413 347 1427 361
rect 1433 347 1447 361
rect 1393 327 1407 341
rect 1453 339 1467 353
rect 1473 347 1487 361
rect 1533 327 1547 341
rect 1553 339 1567 353
rect 1613 347 1627 361
rect 1773 387 1787 401
rect 1753 367 1767 381
rect 1793 367 1807 381
rect 1733 353 1747 367
rect 1813 359 1827 373
rect 1633 339 1647 353
rect 1653 327 1667 341
rect 1673 339 1687 353
rect 1693 327 1707 341
rect 1713 339 1727 353
rect 1753 333 1767 347
rect 1853 339 1867 353
rect 1873 327 1887 341
rect 1893 339 1907 353
rect 1913 347 1927 361
rect 1953 359 1967 373
rect 1973 367 1987 381
rect 2013 373 2027 387
rect 2093 393 2107 407
rect 1993 359 2007 373
rect 2033 359 2047 373
rect 2053 367 2067 381
rect 2033 313 2047 327
rect 2073 359 2087 373
rect 2173 393 2187 407
rect 2113 359 2127 373
rect 2133 367 2147 381
rect 2093 313 2107 327
rect 2153 359 2167 373
rect 2213 347 2227 361
rect 2193 333 2207 347
rect 2253 347 2267 361
rect 2293 359 2307 373
rect 2313 367 2327 381
rect 2233 327 2247 341
rect 2333 359 2347 373
rect 2353 347 2367 361
rect 2453 387 2467 401
rect 2433 367 2447 381
rect 2473 367 2487 381
rect 2393 347 2407 361
rect 2493 359 2507 373
rect 2373 327 2387 341
rect 2653 387 2667 401
rect 2613 359 2627 373
rect 2633 367 2647 381
rect 2673 367 2687 381
rect 2553 339 2567 353
rect 2573 327 2587 341
rect 2693 339 2707 353
rect 2713 327 2727 341
rect 2733 339 2747 353
rect 2753 347 2767 361
rect 2793 347 2807 361
rect 2833 347 2847 361
rect 2893 359 2907 373
rect 2913 367 2927 381
rect 2813 327 2827 341
rect 2933 359 2947 373
rect 2973 367 2987 381
rect 3073 367 3087 381
rect 2993 347 3007 361
rect 3013 339 3027 353
rect 3033 347 3047 361
rect 3093 347 3107 361
rect 3113 339 3127 353
rect 3133 347 3147 361
rect 3173 347 3187 361
rect 3213 347 3227 361
rect 3313 367 3327 381
rect 3193 327 3207 341
rect 3253 339 3267 353
rect 3333 347 3347 361
rect 3273 327 3287 341
rect 3353 339 3367 353
rect 3373 347 3387 361
rect 3413 347 3427 361
rect 3433 339 3447 353
rect 3453 327 3467 341
rect 3473 339 3487 353
rect 3513 347 3527 361
rect 3553 347 3567 361
rect 3593 347 3607 361
rect 3533 327 3547 341
rect 3573 327 3587 341
rect 3673 359 3687 373
rect 3693 367 3707 381
rect 3633 339 3647 353
rect 3713 359 3727 373
rect 3753 359 3767 373
rect 3773 367 3787 381
rect 3793 359 3807 373
rect 3853 367 3867 381
rect 3873 347 3887 361
rect 3893 339 3907 353
rect 3913 347 3927 361
rect 4093 422 4107 436
rect 4233 416 4247 430
rect 3953 339 3967 353
rect 3973 327 3987 341
rect 4013 339 4027 353
rect 4033 327 4047 341
rect 4093 384 4107 398
rect 4073 319 4087 333
rect 4153 347 4167 361
rect 4193 347 4207 361
rect 4093 290 4107 304
rect 4313 359 4327 373
rect 4333 367 4347 381
rect 4353 359 4367 373
rect 4393 367 4407 381
rect 4413 347 4427 361
rect 4433 339 4447 353
rect 4453 347 4467 361
rect 4573 422 4587 436
rect 4713 416 4727 430
rect 4493 339 4507 353
rect 4233 290 4247 304
rect 4513 327 4527 341
rect 4573 384 4587 398
rect 4553 319 4567 333
rect 4633 347 4647 361
rect 4673 347 4687 361
rect 4573 290 4587 304
rect 4713 290 4727 304
rect 113 147 127 161
rect 133 159 147 173
rect 153 147 167 161
rect 33 127 47 141
rect 173 139 187 153
rect 253 139 267 153
rect 273 147 287 161
rect 293 139 307 153
rect 313 139 327 153
rect 333 147 347 161
rect 353 139 367 153
rect 593 173 607 187
rect 53 119 67 133
rect 93 119 107 133
rect 73 99 87 113
rect 233 119 247 133
rect 373 119 387 133
rect 433 127 447 141
rect 453 119 467 133
rect 493 119 507 133
rect 513 119 527 133
rect 553 119 567 133
rect 573 127 587 141
rect 473 99 487 113
rect 533 99 547 113
rect 613 147 627 161
rect 633 159 647 173
rect 653 147 667 161
rect 673 139 687 153
rect 733 139 747 153
rect 753 147 767 161
rect 773 159 787 173
rect 793 147 807 161
rect 813 159 827 173
rect 973 193 987 207
rect 833 147 847 161
rect 593 93 607 107
rect 913 139 927 153
rect 933 147 947 161
rect 953 139 967 153
rect 893 119 907 133
rect 993 147 1007 161
rect 1013 159 1027 173
rect 973 113 987 127
rect 1033 139 1047 153
rect 1053 147 1067 161
rect 1073 139 1087 153
rect 1133 139 1147 153
rect 1153 147 1167 161
rect 1173 139 1187 153
rect 1093 119 1107 133
rect 1193 119 1207 133
rect 1233 119 1247 133
rect 1273 119 1287 133
rect 1293 127 1307 141
rect 1253 99 1267 113
rect 1333 119 1347 133
rect 1373 119 1387 133
rect 1393 127 1407 141
rect 1453 139 1467 153
rect 1473 147 1487 161
rect 1493 159 1507 173
rect 1513 147 1527 161
rect 1353 99 1367 113
rect 1533 119 1547 133
rect 1573 119 1587 133
rect 1593 127 1607 141
rect 1653 139 1667 153
rect 1673 147 1687 161
rect 1693 159 1707 173
rect 1713 147 1727 161
rect 1553 99 1567 113
rect 1733 119 1747 133
rect 1773 119 1787 133
rect 1793 127 1807 141
rect 1833 127 1847 141
rect 1753 99 1767 113
rect 1853 119 1867 133
rect 1873 127 1887 141
rect 1913 139 1927 153
rect 1953 139 1967 153
rect 2013 139 2027 153
rect 2033 127 2047 141
rect 2073 139 2087 153
rect 2093 139 2107 153
rect 2133 139 2147 153
rect 2173 119 2187 133
rect 2213 119 2227 133
rect 2233 127 2247 141
rect 2273 139 2287 153
rect 2293 147 2307 161
rect 2313 139 2327 153
rect 2333 147 2347 161
rect 2353 139 2367 153
rect 2393 139 2407 153
rect 2413 147 2427 161
rect 2433 139 2447 153
rect 2513 139 2527 153
rect 2533 147 2547 161
rect 2553 159 2567 173
rect 2573 147 2587 161
rect 2593 139 2607 153
rect 2613 147 2627 161
rect 2693 159 2707 173
rect 2633 139 2647 153
rect 2713 147 2727 161
rect 2193 99 2207 113
rect 2453 119 2467 133
rect 2653 119 2667 133
rect 2853 159 2867 173
rect 2953 196 2967 210
rect 2873 147 2887 161
rect 2753 119 2767 133
rect 2793 119 2807 133
rect 2813 127 2827 141
rect 2773 99 2787 113
rect 3093 196 3107 210
rect 2993 139 3007 153
rect 3033 139 3047 153
rect 3113 167 3127 181
rect 3093 102 3107 116
rect 3153 159 3167 173
rect 3313 196 3327 210
rect 3173 147 3187 161
rect 3233 147 3247 161
rect 3253 159 3267 173
rect 2953 70 2967 84
rect 3093 64 3107 78
rect 3453 196 3467 210
rect 3353 139 3367 153
rect 3393 139 3407 153
rect 3473 167 3487 181
rect 3453 102 3467 116
rect 3633 196 3647 210
rect 3773 196 3787 210
rect 3553 159 3567 173
rect 3613 167 3627 181
rect 3533 139 3547 153
rect 3573 139 3587 153
rect 3313 70 3327 84
rect 3453 64 3467 78
rect 3633 102 3647 116
rect 3693 139 3707 153
rect 3733 139 3747 153
rect 3833 159 3847 173
rect 3853 147 3867 161
rect 3633 64 3647 78
rect 3773 70 3787 84
rect 3893 139 3907 153
rect 3913 147 3927 161
rect 4013 159 4027 173
rect 4093 159 4107 173
rect 3933 139 3947 153
rect 3993 139 4007 153
rect 3953 119 3967 133
rect 4033 139 4047 153
rect 4073 139 4087 153
rect 4193 159 4207 173
rect 4113 139 4127 153
rect 4173 139 4187 153
rect 4213 139 4227 153
rect 4233 139 4247 153
rect 4253 147 4267 161
rect 4273 139 4287 153
rect 4293 119 4307 133
rect 4353 127 4367 141
rect 4433 147 4447 161
rect 4453 159 4467 173
rect 4493 159 4507 173
rect 4373 119 4387 133
rect 4393 127 4407 141
rect 4473 139 4487 153
rect 4513 139 4527 153
rect 4553 127 4567 141
rect 4653 147 4667 161
rect 4673 159 4687 173
rect 4573 119 4587 133
rect 4593 127 4607 141
rect 4693 127 4707 141
rect 4713 119 4727 133
rect 4733 127 4747 141
<< metal2 >>
rect 3996 4616 4023 4623
rect 36 4487 43 4513
rect 33 4473 47 4487
rect 53 4453 67 4467
rect 56 4407 63 4453
rect 96 4427 103 4453
rect 116 4407 123 4533
rect 176 4487 183 4493
rect 133 4433 147 4447
rect 176 4447 183 4473
rect 196 4467 203 4533
rect 496 4507 503 4513
rect 216 4467 223 4473
rect 193 4453 207 4467
rect 213 4453 227 4467
rect 236 4447 243 4453
rect 136 4367 143 4433
rect 233 4433 247 4447
rect 36 4227 43 4233
rect 33 4213 47 4227
rect 53 4193 67 4207
rect 96 4207 103 4233
rect 156 4227 163 4413
rect 56 4147 63 4193
rect 56 3987 63 4033
rect 76 4027 83 4173
rect 153 4173 167 4187
rect 116 3987 123 4153
rect 156 4107 163 4173
rect 176 4127 183 4393
rect 16 3956 33 3963
rect 16 3703 23 3956
rect 53 3973 67 3987
rect 73 3963 87 3967
rect 93 3963 107 3967
rect 73 3956 107 3963
rect 113 3973 127 3987
rect 73 3953 87 3956
rect 93 3953 107 3956
rect 133 3953 147 3967
rect 56 3727 63 3893
rect 76 3747 83 3953
rect 136 3947 143 3953
rect 136 3747 143 3933
rect 156 3887 163 4073
rect 176 3943 183 4113
rect 196 4067 203 4413
rect 316 4227 323 4453
rect 333 4433 347 4447
rect 376 4447 383 4493
rect 396 4467 403 4473
rect 556 4487 563 4493
rect 656 4487 663 4493
rect 393 4453 407 4467
rect 513 4483 527 4487
rect 496 4476 527 4483
rect 496 4467 503 4476
rect 513 4473 527 4476
rect 533 4453 547 4467
rect 553 4473 567 4487
rect 573 4463 587 4467
rect 573 4456 603 4463
rect 573 4453 587 4456
rect 336 4407 343 4433
rect 416 4287 423 4453
rect 456 4327 463 4453
rect 536 4447 543 4453
rect 507 4436 513 4443
rect 596 4367 603 4456
rect 633 4453 647 4467
rect 653 4473 667 4487
rect 253 4223 267 4227
rect 253 4216 283 4223
rect 253 4213 267 4216
rect 216 3987 223 4013
rect 256 3987 263 4173
rect 276 4087 283 4216
rect 356 4187 363 4273
rect 373 4193 387 4207
rect 296 4147 303 4173
rect 333 4173 347 4187
rect 336 4087 343 4173
rect 376 4127 383 4193
rect 433 4183 447 4187
rect 453 4183 467 4187
rect 433 4176 467 4183
rect 433 4173 447 4176
rect 453 4173 467 4176
rect 436 4107 443 4173
rect 516 4127 523 4193
rect 556 4167 563 4353
rect 576 4207 583 4313
rect 573 4193 587 4207
rect 616 4183 623 4433
rect 636 4427 643 4453
rect 656 4387 663 4433
rect 696 4407 703 4453
rect 716 4443 723 4513
rect 756 4496 863 4503
rect 756 4487 763 4496
rect 856 4487 863 4496
rect 733 4443 747 4447
rect 716 4436 747 4443
rect 776 4447 783 4473
rect 733 4433 747 4436
rect 773 4433 787 4447
rect 836 4447 843 4473
rect 896 4423 903 4533
rect 1056 4516 1143 4523
rect 1056 4507 1063 4516
rect 1136 4507 1143 4516
rect 996 4467 1003 4473
rect 913 4433 927 4447
rect 993 4453 1007 4467
rect 1053 4433 1067 4447
rect 916 4427 923 4433
rect 876 4416 903 4423
rect 656 4207 663 4213
rect 633 4183 647 4187
rect 616 4176 647 4183
rect 653 4193 667 4207
rect 633 4173 647 4176
rect 593 4153 607 4167
rect 716 4167 723 4413
rect 736 4207 743 4373
rect 816 4367 823 4413
rect 833 4223 847 4227
rect 856 4223 863 4413
rect 733 4193 747 4207
rect 813 4193 827 4207
rect 833 4216 863 4223
rect 833 4213 847 4216
rect 596 4147 603 4153
rect 296 4007 303 4053
rect 376 4027 383 4033
rect 373 4013 387 4027
rect 336 4007 343 4013
rect 293 3993 307 4007
rect 213 3973 227 3987
rect 313 3973 327 3987
rect 333 3993 347 4007
rect 416 4007 423 4033
rect 353 3983 367 3987
rect 353 3976 383 3983
rect 353 3973 367 3976
rect 233 3953 247 3967
rect 176 3936 203 3943
rect 33 3703 47 3707
rect 16 3696 47 3703
rect 33 3693 47 3696
rect 36 3627 43 3693
rect 93 3693 107 3707
rect 133 3693 147 3707
rect 76 3667 83 3693
rect 96 3647 103 3693
rect 56 3507 63 3633
rect 116 3627 123 3673
rect 136 3667 143 3693
rect 33 3473 47 3487
rect 53 3493 67 3507
rect 16 3427 23 3473
rect 16 3207 23 3393
rect 36 3287 43 3473
rect 96 3463 103 3613
rect 116 3487 123 3593
rect 76 3456 103 3463
rect 36 3183 43 3273
rect 56 3184 64 3296
rect 16 3176 43 3183
rect 16 2947 23 3176
rect 76 3047 83 3456
rect 96 3267 103 3433
rect 116 3267 123 3473
rect 136 3444 144 3556
rect 96 3167 103 3193
rect 116 3123 123 3253
rect 133 3213 147 3227
rect 136 3207 143 3213
rect 156 3187 163 3693
rect 176 3667 183 3873
rect 176 3527 183 3533
rect 173 3513 187 3527
rect 196 3483 203 3936
rect 236 3903 243 3953
rect 256 3903 263 3913
rect 316 3907 323 3973
rect 236 3896 263 3903
rect 256 3703 263 3896
rect 356 3727 363 3953
rect 376 3887 383 3976
rect 393 3973 407 3987
rect 413 3993 427 4007
rect 473 4003 487 4007
rect 456 3996 487 4003
rect 396 3907 403 3973
rect 436 3927 443 3993
rect 456 3947 463 3996
rect 473 3993 487 3996
rect 533 3953 547 3967
rect 573 3953 587 3967
rect 536 3927 543 3953
rect 576 3947 583 3953
rect 596 3907 603 4113
rect 656 4007 663 4053
rect 653 3993 667 4007
rect 273 3703 287 3707
rect 256 3696 287 3703
rect 273 3693 287 3696
rect 373 3693 387 3707
rect 236 3647 243 3673
rect 213 3523 227 3527
rect 213 3516 243 3523
rect 213 3513 227 3516
rect 176 3476 203 3483
rect 176 3247 183 3476
rect 195 3278 203 3302
rect 136 3147 143 3173
rect 176 3143 183 3213
rect 195 3184 203 3264
rect 236 3207 243 3516
rect 256 3367 263 3673
rect 275 3476 283 3556
rect 293 3513 307 3527
rect 275 3438 283 3462
rect 296 3447 303 3513
rect 296 3407 303 3433
rect 176 3136 203 3143
rect 116 3116 143 3123
rect 53 3013 67 3027
rect 73 3033 87 3047
rect 16 2707 23 2773
rect 36 2767 43 2993
rect 56 2987 63 3013
rect 136 3003 143 3116
rect 156 3047 163 3053
rect 153 3033 167 3047
rect 136 2996 163 3003
rect 56 2767 63 2913
rect 76 2847 83 2993
rect 96 2823 103 2973
rect 76 2816 103 2823
rect 53 2713 67 2727
rect 36 2587 43 2713
rect 56 2707 63 2713
rect 16 2547 23 2553
rect 13 2533 27 2547
rect 36 2527 43 2573
rect 56 2547 63 2653
rect 76 2567 83 2816
rect 156 2787 163 2996
rect 173 2993 187 3007
rect 176 2947 183 2993
rect 176 2843 183 2933
rect 196 2867 203 3136
rect 213 3043 227 3047
rect 236 3043 243 3113
rect 256 3087 263 3333
rect 316 3327 323 3633
rect 356 3587 363 3693
rect 376 3667 383 3693
rect 416 3687 423 3753
rect 473 3743 487 3747
rect 456 3736 487 3743
rect 433 3693 447 3707
rect 436 3647 443 3693
rect 456 3647 463 3736
rect 473 3733 487 3736
rect 536 3707 543 3893
rect 556 3747 563 3753
rect 596 3747 603 3753
rect 553 3733 567 3747
rect 593 3733 607 3747
rect 636 3727 643 3753
rect 633 3713 647 3727
rect 516 3667 523 3693
rect 336 3503 343 3573
rect 376 3547 383 3613
rect 536 3587 543 3673
rect 373 3543 387 3547
rect 373 3536 403 3543
rect 373 3533 387 3536
rect 353 3503 367 3507
rect 336 3496 367 3503
rect 353 3493 367 3496
rect 376 3467 383 3493
rect 396 3343 403 3536
rect 516 3527 523 3533
rect 513 3513 527 3527
rect 413 3473 427 3487
rect 453 3483 467 3487
rect 476 3483 483 3513
rect 453 3476 483 3483
rect 453 3473 467 3476
rect 416 3467 423 3473
rect 376 3336 403 3343
rect 296 3247 303 3273
rect 336 3247 343 3273
rect 376 3247 383 3336
rect 456 3327 463 3473
rect 396 3307 403 3313
rect 396 3267 403 3273
rect 393 3253 407 3267
rect 273 3213 287 3227
rect 293 3233 307 3247
rect 313 3213 327 3227
rect 333 3233 347 3247
rect 276 3127 283 3213
rect 316 3203 323 3213
rect 316 3196 343 3203
rect 336 3187 343 3196
rect 213 3036 243 3043
rect 213 3033 227 3036
rect 176 2836 203 2843
rect 136 2767 143 2773
rect 196 2767 203 2836
rect 216 2787 223 2993
rect 236 2827 243 3036
rect 253 3033 267 3047
rect 256 2907 263 3033
rect 277 2996 285 3076
rect 296 3027 303 3133
rect 277 2958 285 2982
rect 93 2753 107 2767
rect 96 2667 103 2753
rect 133 2753 147 2767
rect 153 2733 167 2747
rect 213 2733 227 2747
rect 276 2747 283 2813
rect 296 2787 303 2993
rect 316 2927 323 3173
rect 333 3043 347 3047
rect 356 3043 363 3193
rect 376 3187 383 3213
rect 333 3036 363 3043
rect 333 3033 347 3036
rect 356 2887 363 3036
rect 376 2967 383 2993
rect 396 2943 403 3153
rect 436 3127 443 3213
rect 456 3187 463 3293
rect 497 3278 505 3302
rect 476 3227 483 3253
rect 497 3184 505 3264
rect 416 2964 424 3076
rect 436 2967 443 3113
rect 376 2936 403 2943
rect 336 2787 343 2793
rect 376 2787 383 2936
rect 313 2753 327 2767
rect 333 2773 347 2787
rect 413 2783 427 2787
rect 396 2776 427 2783
rect 33 2513 47 2527
rect 73 2513 87 2527
rect 16 2327 23 2493
rect 36 2327 43 2393
rect 76 2343 83 2513
rect 96 2363 103 2613
rect 156 2607 163 2733
rect 176 2627 183 2733
rect 196 2683 203 2713
rect 216 2707 223 2733
rect 196 2676 223 2683
rect 173 2563 187 2567
rect 173 2556 203 2563
rect 173 2553 187 2556
rect 96 2356 123 2363
rect 76 2336 103 2343
rect 96 2327 103 2336
rect 33 2303 47 2307
rect 16 2296 47 2303
rect 16 2187 23 2296
rect 33 2293 47 2296
rect 73 2293 87 2307
rect 76 2267 83 2293
rect 56 2256 73 2263
rect 16 2007 23 2173
rect 36 2087 43 2253
rect 56 2107 63 2256
rect 76 2087 83 2093
rect 33 2073 47 2087
rect 73 2073 87 2087
rect 16 1727 23 1873
rect 36 1823 43 1853
rect 56 1847 63 2073
rect 96 2063 103 2253
rect 116 2087 123 2356
rect 136 2347 143 2353
rect 196 2307 203 2556
rect 216 2407 223 2676
rect 256 2587 263 2593
rect 253 2573 267 2587
rect 296 2567 303 2713
rect 316 2667 323 2753
rect 356 2727 363 2773
rect 396 2767 403 2776
rect 413 2773 427 2776
rect 396 2723 403 2753
rect 376 2716 403 2723
rect 293 2563 307 2567
rect 276 2556 307 2563
rect 256 2303 263 2533
rect 276 2367 283 2556
rect 293 2553 307 2556
rect 336 2467 343 2693
rect 356 2567 363 2613
rect 353 2553 367 2567
rect 376 2527 383 2716
rect 416 2667 423 2733
rect 436 2587 443 2613
rect 456 2587 463 3153
rect 476 3047 483 3093
rect 516 3087 523 3313
rect 536 3067 543 3353
rect 556 3307 563 3473
rect 553 3213 567 3227
rect 556 3207 563 3213
rect 576 3167 583 3693
rect 613 3673 627 3687
rect 656 3683 663 3933
rect 696 3927 703 4153
rect 776 4147 783 4193
rect 816 4187 823 4193
rect 856 4187 863 4216
rect 876 4167 883 4416
rect 956 4367 963 4433
rect 1056 4407 1063 4433
rect 1076 4367 1083 4493
rect 1133 4453 1147 4467
rect 1096 4427 1103 4453
rect 1136 4447 1143 4453
rect 1176 4427 1183 4473
rect 1236 4467 1243 4553
rect 1276 4467 1283 4493
rect 1296 4487 1303 4533
rect 1293 4473 1307 4487
rect 916 4227 923 4353
rect 1013 4223 1027 4227
rect 996 4216 1027 4223
rect 916 4207 923 4213
rect 913 4193 927 4207
rect 933 4173 947 4187
rect 973 4183 987 4187
rect 996 4183 1003 4216
rect 1013 4213 1027 4216
rect 1156 4227 1163 4353
rect 1033 4193 1047 4207
rect 973 4176 1003 4183
rect 973 4173 987 4176
rect 936 4167 943 4173
rect 1036 4147 1043 4193
rect 716 3963 723 4013
rect 776 4007 783 4133
rect 796 3987 803 4053
rect 856 3987 863 4033
rect 733 3963 747 3967
rect 716 3956 747 3963
rect 793 3973 807 3987
rect 733 3953 747 3956
rect 853 3973 867 3987
rect 873 3963 887 3967
rect 896 3963 903 4133
rect 936 3987 943 4033
rect 956 4007 963 4033
rect 1056 4007 1063 4213
rect 1073 4193 1087 4207
rect 1093 4203 1107 4207
rect 1093 4196 1123 4203
rect 1093 4193 1107 4196
rect 1076 4127 1083 4193
rect 953 3993 967 4007
rect 873 3956 903 3963
rect 933 3973 947 3987
rect 1053 3993 1067 4007
rect 1076 3987 1083 4053
rect 1073 3973 1087 3987
rect 873 3953 887 3956
rect 756 3767 763 3933
rect 773 3743 787 3747
rect 756 3736 787 3743
rect 813 3743 827 3747
rect 836 3743 843 3773
rect 756 3707 763 3736
rect 773 3733 787 3736
rect 813 3736 843 3743
rect 813 3733 827 3736
rect 713 3703 727 3707
rect 713 3696 733 3703
rect 713 3693 727 3696
rect 836 3687 843 3736
rect 656 3676 683 3683
rect 596 3507 603 3573
rect 616 3527 623 3673
rect 656 3527 663 3593
rect 676 3567 683 3676
rect 696 3627 703 3673
rect 613 3513 627 3527
rect 593 3493 607 3507
rect 633 3493 647 3507
rect 596 3267 603 3293
rect 596 3107 603 3173
rect 616 3167 623 3393
rect 636 3347 643 3493
rect 673 3473 687 3487
rect 713 3473 727 3487
rect 676 3467 683 3473
rect 636 3184 644 3296
rect 656 3187 663 3253
rect 473 3033 487 3047
rect 493 3013 507 3027
rect 433 2573 447 2587
rect 453 2533 467 2547
rect 316 2327 323 2353
rect 356 2327 363 2513
rect 416 2347 423 2413
rect 236 2296 263 2303
rect 236 2287 243 2296
rect 133 2273 147 2287
rect 136 2267 143 2273
rect 153 2253 167 2267
rect 193 2253 207 2267
rect 213 2253 227 2267
rect 253 2253 267 2267
rect 156 2207 163 2253
rect 196 2247 203 2253
rect 216 2247 223 2253
rect 176 2087 183 2133
rect 216 2087 223 2213
rect 236 2087 243 2213
rect 256 2087 263 2253
rect 276 2227 283 2273
rect 296 2247 303 2293
rect 333 2293 347 2307
rect 373 2303 387 2307
rect 336 2267 343 2293
rect 373 2296 403 2303
rect 373 2293 387 2296
rect 336 2247 343 2253
rect 113 2063 127 2067
rect 96 2056 127 2063
rect 113 2053 127 2056
rect 153 2053 167 2067
rect 233 2063 247 2067
rect 256 2063 263 2073
rect 276 2067 283 2153
rect 316 2107 323 2173
rect 356 2107 363 2193
rect 313 2093 327 2107
rect 76 1827 83 2033
rect 96 1887 103 2033
rect 116 1847 123 1993
rect 36 1816 63 1823
rect 56 1807 63 1816
rect 96 1807 103 1813
rect 156 1807 163 2053
rect 213 2033 227 2047
rect 233 2056 263 2063
rect 233 2053 247 2056
rect 333 2053 347 2067
rect 176 1987 183 2033
rect 216 1967 223 2033
rect 236 1947 243 2013
rect 216 1847 223 1853
rect 236 1847 243 1913
rect 296 1883 303 1933
rect 316 1907 323 2053
rect 336 2047 343 2053
rect 296 1876 323 1883
rect 236 1827 243 1833
rect 233 1813 247 1827
rect 273 1823 287 1827
rect 296 1823 303 1853
rect 33 1773 47 1787
rect 53 1793 67 1807
rect 93 1793 107 1807
rect 113 1773 127 1787
rect 133 1773 147 1787
rect 173 1773 187 1787
rect 36 1747 43 1773
rect 96 1627 103 1753
rect 116 1707 123 1773
rect 136 1727 143 1773
rect 176 1747 183 1773
rect 136 1687 143 1713
rect 176 1627 183 1733
rect 53 1623 67 1627
rect 53 1616 83 1623
rect 53 1613 67 1616
rect 16 1147 23 1593
rect 76 1407 83 1616
rect 176 1587 183 1613
rect 173 1573 187 1587
rect 116 1567 123 1573
rect 56 1347 63 1393
rect 136 1387 143 1573
rect 196 1567 203 1773
rect 216 1747 223 1813
rect 273 1816 303 1823
rect 273 1813 287 1816
rect 256 1767 263 1793
rect 276 1707 283 1773
rect 233 1553 247 1567
rect 256 1563 263 1693
rect 276 1627 283 1633
rect 296 1627 303 1816
rect 316 1727 323 1876
rect 376 1867 383 2253
rect 396 2227 403 2296
rect 416 2287 423 2333
rect 436 2287 443 2533
rect 456 2527 463 2533
rect 476 2487 483 2973
rect 496 2947 503 3013
rect 536 2807 543 2953
rect 556 2927 563 3093
rect 576 3067 583 3093
rect 596 3047 603 3073
rect 613 2993 627 3007
rect 616 2947 623 2993
rect 556 2827 563 2833
rect 556 2783 563 2813
rect 576 2787 583 2893
rect 636 2883 643 3133
rect 656 2907 663 3153
rect 676 3147 683 3353
rect 696 3243 703 3453
rect 716 3387 723 3473
rect 736 3367 743 3553
rect 756 3547 763 3613
rect 756 3527 763 3533
rect 796 3527 803 3633
rect 836 3527 843 3533
rect 753 3513 767 3527
rect 773 3493 787 3507
rect 793 3513 807 3527
rect 813 3493 827 3507
rect 756 3247 763 3373
rect 776 3347 783 3493
rect 816 3447 823 3493
rect 713 3243 727 3247
rect 696 3236 727 3243
rect 713 3233 727 3236
rect 753 3233 767 3247
rect 773 3213 787 3227
rect 776 3203 783 3213
rect 796 3207 803 3273
rect 816 3267 823 3433
rect 856 3407 863 3913
rect 876 3807 883 3933
rect 876 3747 883 3793
rect 873 3733 887 3747
rect 893 3723 907 3727
rect 956 3727 963 3773
rect 976 3727 983 3953
rect 1036 3947 1043 3973
rect 1096 3967 1103 4173
rect 1116 3907 1123 4196
rect 1133 4193 1147 4207
rect 1153 4213 1167 4227
rect 1196 4223 1203 4453
rect 1213 4433 1227 4447
rect 1233 4453 1247 4467
rect 1216 4387 1223 4433
rect 1256 4407 1263 4433
rect 1356 4427 1363 4493
rect 1436 4487 1443 4513
rect 1456 4507 1463 4533
rect 1413 4453 1427 4467
rect 1433 4473 1447 4487
rect 1416 4407 1423 4453
rect 1456 4443 1463 4493
rect 1536 4487 1543 4553
rect 1533 4473 1547 4487
rect 1496 4467 1503 4473
rect 1473 4443 1487 4447
rect 1456 4436 1487 4443
rect 1493 4453 1507 4467
rect 1616 4467 1623 4513
rect 1613 4453 1627 4467
rect 1473 4433 1487 4436
rect 1556 4407 1563 4453
rect 1596 4427 1603 4453
rect 1636 4447 1643 4533
rect 1633 4433 1647 4447
rect 1696 4447 1703 4513
rect 1816 4507 1823 4513
rect 1956 4507 1963 4513
rect 1733 4483 1747 4487
rect 1716 4476 1747 4483
rect 1673 4433 1687 4447
rect 1676 4267 1683 4433
rect 1396 4227 1403 4233
rect 1213 4223 1227 4227
rect 1196 4216 1227 4223
rect 1253 4223 1267 4227
rect 1136 4147 1143 4193
rect 1196 4147 1203 4216
rect 1213 4213 1227 4216
rect 1253 4216 1283 4223
rect 1253 4213 1267 4216
rect 1276 4187 1283 4216
rect 1333 4213 1347 4227
rect 1336 4187 1343 4213
rect 1353 4193 1367 4207
rect 1393 4213 1407 4227
rect 1413 4193 1427 4207
rect 1513 4223 1527 4227
rect 1153 4023 1167 4027
rect 1153 4016 1183 4023
rect 1153 4013 1167 4016
rect 1176 3807 1183 4016
rect 1216 3987 1223 4033
rect 1236 4027 1243 4173
rect 1273 4023 1287 4027
rect 1256 4016 1287 4023
rect 1213 3973 1227 3987
rect 1236 3967 1243 4013
rect 1256 3987 1263 4016
rect 1273 4013 1287 4016
rect 1336 3987 1343 4113
rect 1356 4107 1363 4193
rect 1253 3983 1267 3987
rect 1253 3976 1283 3983
rect 1253 3973 1267 3976
rect 1233 3953 1247 3967
rect 1276 3907 1283 3976
rect 1356 3967 1363 4013
rect 1376 3987 1383 4033
rect 1396 4007 1403 4173
rect 1416 4127 1423 4193
rect 1373 3973 1387 3987
rect 1353 3953 1367 3967
rect 1416 3947 1423 4093
rect 1436 3987 1443 4013
rect 1433 3973 1447 3987
rect 1456 3967 1463 4133
rect 1476 4027 1483 4213
rect 1493 4193 1507 4207
rect 1513 4216 1543 4223
rect 1513 4213 1527 4216
rect 1496 4167 1503 4193
rect 1536 4087 1543 4216
rect 1556 4207 1563 4233
rect 1716 4223 1723 4476
rect 1733 4473 1747 4476
rect 1813 4493 1827 4507
rect 1753 4453 1767 4467
rect 1793 4453 1807 4467
rect 1833 4453 1847 4467
rect 1953 4493 1967 4507
rect 1933 4453 1947 4467
rect 1973 4453 1987 4467
rect 2016 4483 2023 4513
rect 2056 4507 2063 4513
rect 2053 4493 2067 4507
rect 2113 4503 2127 4507
rect 2033 4483 2047 4487
rect 2016 4476 2047 4483
rect 2096 4496 2127 4503
rect 2073 4483 2087 4487
rect 2096 4483 2103 4496
rect 2016 4467 2023 4476
rect 2033 4473 2047 4476
rect 2073 4476 2103 4483
rect 2113 4493 2127 4496
rect 2176 4487 2183 4493
rect 2073 4473 2087 4476
rect 1756 4407 1763 4453
rect 1796 4327 1803 4453
rect 1836 4447 1843 4453
rect 1936 4327 1943 4453
rect 1976 4447 1983 4453
rect 1716 4216 1743 4223
rect 1736 4207 1743 4216
rect 1556 4183 1563 4193
rect 1573 4183 1587 4187
rect 1556 4176 1587 4183
rect 1573 4173 1587 4176
rect 1613 4173 1627 4187
rect 1653 4173 1667 4187
rect 1593 4153 1607 4167
rect 1496 4016 1563 4023
rect 1496 4003 1503 4016
rect 1476 3996 1503 4003
rect 1476 3987 1483 3996
rect 1473 3973 1487 3987
rect 996 3727 1003 3753
rect 1036 3747 1043 3793
rect 893 3716 923 3723
rect 893 3713 907 3716
rect 916 3687 923 3716
rect 933 3713 947 3727
rect 953 3713 967 3727
rect 993 3713 1007 3727
rect 936 3707 943 3713
rect 936 3687 943 3693
rect 1056 3707 1063 3713
rect 1076 3687 1083 3733
rect 1153 3723 1167 3727
rect 1136 3716 1167 3723
rect 836 3247 843 3293
rect 876 3267 883 3493
rect 916 3367 923 3673
rect 936 3483 943 3653
rect 976 3567 983 3673
rect 1076 3607 1083 3633
rect 1096 3607 1103 3713
rect 1136 3707 1143 3716
rect 1153 3713 1167 3716
rect 1213 3693 1227 3707
rect 1216 3687 1223 3693
rect 956 3523 963 3553
rect 996 3527 1003 3573
rect 956 3516 983 3523
rect 976 3507 983 3516
rect 1016 3507 1023 3533
rect 1096 3527 1103 3533
rect 953 3483 967 3487
rect 936 3476 967 3483
rect 973 3493 987 3507
rect 1073 3493 1087 3507
rect 1093 3513 1107 3527
rect 1116 3507 1123 3573
rect 1136 3527 1143 3613
rect 1156 3547 1163 3573
rect 1236 3547 1243 3893
rect 1336 3747 1343 3853
rect 1333 3733 1347 3747
rect 1393 3713 1407 3727
rect 1396 3687 1403 3713
rect 1416 3687 1423 3753
rect 1476 3707 1483 3933
rect 1516 3867 1523 3993
rect 1556 3987 1563 4016
rect 1596 4007 1603 4153
rect 1616 4107 1623 4173
rect 1656 4107 1663 4173
rect 1693 4173 1707 4187
rect 1713 4173 1727 4187
rect 1773 4203 1787 4207
rect 1796 4203 1803 4233
rect 1773 4196 1803 4203
rect 1773 4193 1787 4196
rect 1853 4193 1867 4207
rect 1896 4207 1903 4313
rect 1916 4207 1923 4213
rect 1913 4193 1927 4207
rect 1936 4203 1943 4233
rect 1953 4203 1967 4207
rect 1936 4196 1967 4203
rect 1953 4193 1967 4196
rect 1993 4193 2007 4207
rect 1696 4007 1703 4173
rect 1716 4127 1723 4173
rect 1716 4007 1723 4093
rect 1816 4067 1823 4193
rect 1856 4147 1863 4193
rect 1533 3953 1547 3967
rect 1553 3973 1567 3987
rect 1713 3993 1727 4007
rect 1573 3953 1587 3967
rect 1733 3963 1747 3967
rect 1716 3956 1747 3963
rect 1536 3947 1543 3953
rect 1576 3867 1583 3953
rect 1256 3667 1263 3673
rect 1153 3533 1167 3547
rect 1133 3513 1147 3527
rect 1173 3523 1187 3527
rect 1173 3516 1203 3523
rect 1173 3513 1187 3516
rect 953 3473 967 3476
rect 1036 3487 1043 3493
rect 936 3407 943 3453
rect 1076 3447 1083 3493
rect 916 3267 923 3273
rect 913 3253 927 3267
rect 813 3213 827 3227
rect 833 3233 847 3247
rect 816 3207 823 3213
rect 756 3196 783 3203
rect 636 2876 663 2883
rect 616 2787 623 2833
rect 536 2776 563 2783
rect 536 2767 543 2776
rect 496 2747 503 2753
rect 513 2733 527 2747
rect 533 2753 547 2767
rect 593 2753 607 2767
rect 613 2773 627 2787
rect 516 2603 523 2733
rect 507 2596 523 2603
rect 516 2547 523 2573
rect 536 2567 543 2713
rect 536 2547 543 2553
rect 556 2547 563 2593
rect 493 2513 507 2527
rect 513 2533 527 2547
rect 553 2533 567 2547
rect 496 2427 503 2513
rect 576 2507 583 2733
rect 596 2607 603 2753
rect 616 2707 623 2733
rect 656 2707 663 2876
rect 676 2827 683 2973
rect 696 2767 703 2953
rect 716 2807 723 2953
rect 736 2847 743 3193
rect 756 3167 763 3196
rect 776 3067 783 3173
rect 773 3053 787 3067
rect 796 3047 803 3093
rect 836 3083 843 3193
rect 876 3167 883 3173
rect 836 3076 863 3083
rect 836 3047 843 3053
rect 856 3047 863 3076
rect 793 3033 807 3047
rect 836 3027 843 3033
rect 833 3013 847 3027
rect 853 2993 867 3007
rect 736 2783 743 2833
rect 756 2807 763 2933
rect 776 2787 783 2973
rect 856 2847 863 2993
rect 876 2967 883 3153
rect 896 2987 903 3213
rect 976 3167 983 3353
rect 996 3247 1003 3273
rect 1016 3267 1023 3393
rect 1096 3387 1103 3473
rect 1096 3347 1103 3373
rect 1013 3253 1027 3267
rect 1033 3243 1047 3247
rect 1033 3236 1063 3243
rect 1033 3233 1047 3236
rect 1056 3223 1063 3236
rect 1056 3216 1073 3223
rect 916 3027 923 3113
rect 936 3047 943 3153
rect 933 3033 947 3047
rect 913 3013 927 3027
rect 953 3013 967 3027
rect 773 2783 787 2787
rect 716 2776 743 2783
rect 756 2776 787 2783
rect 693 2753 707 2767
rect 676 2683 683 2733
rect 656 2676 683 2683
rect 616 2587 623 2613
rect 616 2567 623 2573
rect 656 2567 663 2676
rect 716 2587 723 2776
rect 756 2767 763 2776
rect 773 2773 787 2776
rect 753 2753 767 2767
rect 793 2753 807 2767
rect 836 2767 843 2813
rect 613 2553 627 2567
rect 596 2547 603 2553
rect 593 2533 607 2547
rect 633 2533 647 2547
rect 653 2553 667 2567
rect 693 2563 707 2567
rect 676 2556 707 2563
rect 576 2427 583 2493
rect 456 2287 463 2353
rect 516 2303 523 2313
rect 496 2296 523 2303
rect 413 2273 427 2287
rect 453 2273 467 2287
rect 396 2103 403 2213
rect 413 2103 427 2107
rect 396 2096 427 2103
rect 413 2093 427 2096
rect 456 2087 463 2113
rect 476 2107 483 2233
rect 453 2073 467 2087
rect 496 2083 503 2296
rect 513 2253 527 2267
rect 573 2273 587 2287
rect 516 2243 523 2253
rect 516 2236 543 2243
rect 476 2076 503 2083
rect 396 1887 403 2033
rect 416 1847 423 2053
rect 436 2047 443 2053
rect 353 1793 367 1807
rect 456 1823 463 1853
rect 476 1847 483 2076
rect 493 2063 507 2067
rect 516 2063 523 2213
rect 536 2167 543 2236
rect 576 2227 583 2273
rect 596 2267 603 2473
rect 616 2263 623 2513
rect 636 2327 643 2533
rect 676 2387 683 2556
rect 693 2553 707 2556
rect 776 2547 783 2693
rect 796 2647 803 2753
rect 816 2667 823 2733
rect 796 2587 803 2613
rect 713 2533 727 2547
rect 696 2363 703 2513
rect 716 2487 723 2533
rect 773 2533 787 2547
rect 793 2513 807 2527
rect 756 2407 763 2513
rect 796 2507 803 2513
rect 816 2487 823 2653
rect 836 2567 843 2653
rect 856 2547 863 2613
rect 876 2547 883 2893
rect 896 2787 903 2833
rect 893 2773 907 2787
rect 896 2567 903 2733
rect 936 2647 943 2993
rect 956 2947 963 3013
rect 996 3007 1003 3093
rect 1016 3027 1023 3053
rect 1036 3047 1043 3073
rect 1076 3047 1083 3093
rect 1033 3033 1047 3047
rect 1013 3013 1027 3027
rect 1053 3013 1067 3027
rect 1073 3033 1087 3047
rect 1096 3043 1103 3333
rect 1136 3307 1143 3333
rect 1136 3267 1143 3293
rect 1133 3253 1147 3267
rect 1116 3047 1123 3133
rect 1136 3067 1143 3153
rect 1156 3067 1163 3493
rect 1196 3487 1203 3516
rect 1213 3473 1227 3487
rect 1216 3407 1223 3473
rect 1256 3427 1263 3473
rect 1216 3327 1223 3393
rect 1176 3267 1183 3293
rect 1276 3267 1283 3553
rect 1376 3527 1383 3633
rect 1373 3513 1387 3527
rect 1393 3493 1407 3507
rect 1396 3483 1403 3493
rect 1387 3476 1403 3483
rect 1376 3367 1383 3473
rect 1213 3253 1227 3267
rect 1193 3233 1207 3247
rect 1173 3213 1187 3227
rect 1176 3207 1183 3213
rect 1176 3107 1183 3193
rect 1196 3087 1203 3233
rect 1216 3167 1223 3253
rect 1233 3233 1247 3247
rect 1236 3167 1243 3233
rect 1133 3053 1147 3067
rect 1113 3043 1127 3047
rect 1096 3036 1127 3043
rect 1153 3043 1167 3047
rect 1176 3043 1183 3053
rect 1056 2967 1063 3013
rect 853 2533 867 2547
rect 893 2543 907 2547
rect 916 2543 923 2573
rect 936 2547 943 2633
rect 956 2607 963 2773
rect 1016 2767 1023 2953
rect 1096 2947 1103 3036
rect 1113 3033 1127 3036
rect 1153 3036 1183 3043
rect 1153 3033 1167 3036
rect 1176 3027 1183 3036
rect 1196 3027 1203 3073
rect 1216 3047 1223 3113
rect 1256 3047 1263 3073
rect 1276 3047 1283 3233
rect 1293 3213 1307 3227
rect 1333 3213 1347 3227
rect 1296 3087 1303 3213
rect 1336 3207 1343 3213
rect 1376 3123 1383 3353
rect 1436 3267 1443 3333
rect 1413 3233 1427 3247
rect 1433 3253 1447 3267
rect 1416 3167 1423 3233
rect 1356 3116 1383 3123
rect 1213 3033 1227 3047
rect 1193 3013 1207 3027
rect 1253 3033 1267 3047
rect 1296 3027 1303 3073
rect 1176 2887 1183 3013
rect 1293 3013 1307 3027
rect 1313 2993 1327 3007
rect 1356 3003 1363 3116
rect 1396 3103 1403 3133
rect 1376 3096 1403 3103
rect 1376 3047 1383 3096
rect 1373 3033 1387 3047
rect 1436 3027 1443 3213
rect 1456 3207 1463 3673
rect 1556 3667 1563 3693
rect 1576 3687 1583 3733
rect 1636 3727 1643 3753
rect 1633 3713 1647 3727
rect 1716 3707 1723 3956
rect 1733 3953 1747 3956
rect 1756 3727 1763 3993
rect 1516 3444 1524 3556
rect 1536 3463 1543 3593
rect 1536 3456 1563 3463
rect 1476 3167 1483 3393
rect 1496 3247 1503 3253
rect 1493 3233 1507 3247
rect 1516 3187 1523 3253
rect 1556 3247 1563 3456
rect 1496 3107 1503 3173
rect 1393 3013 1407 3027
rect 1356 2996 1383 3003
rect 1056 2787 1063 2813
rect 1053 2773 1067 2787
rect 973 2753 987 2767
rect 976 2747 983 2753
rect 993 2733 1007 2747
rect 1073 2753 1087 2767
rect 1076 2747 1083 2753
rect 1033 2733 1047 2747
rect 976 2587 983 2653
rect 996 2647 1003 2733
rect 956 2567 963 2573
rect 1016 2567 1023 2713
rect 1036 2707 1043 2733
rect 953 2553 967 2567
rect 893 2536 923 2543
rect 893 2533 907 2536
rect 933 2533 947 2547
rect 973 2533 987 2547
rect 1036 2547 1043 2613
rect 1056 2567 1063 2733
rect 1116 2707 1123 2873
rect 1136 2687 1143 2813
rect 1196 2787 1203 2793
rect 1196 2767 1203 2773
rect 1153 2753 1167 2767
rect 1156 2747 1163 2753
rect 1193 2753 1207 2767
rect 1213 2733 1227 2747
rect 1236 2743 1243 2973
rect 1256 2787 1263 2993
rect 1277 2798 1285 2822
rect 1253 2743 1267 2747
rect 1236 2736 1267 2743
rect 1216 2707 1223 2733
rect 1096 2607 1103 2653
rect 1236 2647 1243 2736
rect 1253 2733 1267 2736
rect 1277 2704 1285 2784
rect 1296 2727 1303 2953
rect 1316 2827 1323 2993
rect 676 2356 703 2363
rect 656 2287 663 2293
rect 676 2287 683 2356
rect 736 2287 743 2293
rect 633 2263 647 2267
rect 616 2256 647 2263
rect 653 2273 667 2287
rect 633 2253 647 2256
rect 733 2273 747 2287
rect 673 2243 687 2247
rect 656 2236 687 2243
rect 556 2083 563 2193
rect 576 2187 583 2213
rect 656 2207 663 2236
rect 673 2233 687 2236
rect 713 2233 727 2247
rect 616 2136 663 2143
rect 536 2076 563 2083
rect 536 2067 543 2076
rect 493 2056 523 2063
rect 493 2053 507 2056
rect 533 2053 547 2067
rect 456 1816 483 1823
rect 436 1807 443 1813
rect 476 1807 483 1816
rect 393 1793 407 1807
rect 273 1563 287 1567
rect 256 1556 287 1563
rect 56 1327 63 1333
rect 96 1327 103 1373
rect 196 1367 203 1453
rect 236 1387 243 1553
rect 256 1367 263 1556
rect 273 1553 287 1556
rect 313 1553 327 1567
rect 316 1547 323 1553
rect 276 1367 283 1533
rect 296 1367 303 1433
rect 336 1363 343 1773
rect 356 1767 363 1793
rect 396 1783 403 1793
rect 413 1783 427 1787
rect 396 1776 427 1783
rect 433 1793 447 1807
rect 413 1773 427 1776
rect 473 1793 487 1807
rect 356 1427 363 1653
rect 376 1607 383 1773
rect 416 1747 423 1773
rect 516 1747 523 1993
rect 556 1783 563 1913
rect 576 1867 583 2113
rect 616 2047 623 2136
rect 636 2067 643 2113
rect 656 2087 663 2136
rect 613 2033 627 2047
rect 653 2033 667 2047
rect 547 1776 563 1783
rect 616 1787 623 1893
rect 593 1773 607 1787
rect 596 1767 603 1773
rect 636 1767 643 2013
rect 656 1987 663 2033
rect 676 1927 683 2213
rect 716 2187 723 2233
rect 756 2147 763 2353
rect 716 2107 723 2113
rect 776 2107 783 2453
rect 816 2307 823 2393
rect 813 2293 827 2307
rect 796 2127 803 2253
rect 836 2247 843 2473
rect 876 2307 883 2393
rect 916 2307 923 2453
rect 873 2293 887 2307
rect 893 2273 907 2287
rect 713 2093 727 2107
rect 753 2083 767 2087
rect 733 2053 747 2067
rect 753 2076 783 2083
rect 753 2073 767 2076
rect 696 1967 703 2053
rect 716 1907 723 2033
rect 736 2007 743 2053
rect 676 1807 683 1813
rect 653 1773 667 1787
rect 396 1607 403 1713
rect 416 1647 423 1733
rect 393 1593 407 1607
rect 356 1367 363 1393
rect 316 1356 343 1363
rect 133 1333 147 1347
rect 33 1293 47 1307
rect 53 1313 67 1327
rect 36 1127 43 1293
rect 136 1287 143 1333
rect 153 1313 167 1327
rect 273 1343 287 1347
rect 213 1323 227 1327
rect 196 1316 227 1323
rect 156 1307 163 1313
rect 56 1127 63 1253
rect 96 1127 103 1133
rect 116 1127 123 1133
rect 156 1127 163 1153
rect 176 1127 183 1293
rect 53 1113 67 1127
rect 16 947 23 1113
rect 93 1113 107 1127
rect 113 1113 127 1127
rect 153 1113 167 1127
rect 173 1103 187 1107
rect 196 1103 203 1316
rect 213 1313 227 1316
rect 216 1187 223 1293
rect 236 1147 243 1333
rect 273 1336 303 1343
rect 273 1333 287 1336
rect 216 1107 223 1113
rect 173 1096 203 1103
rect 173 1093 187 1096
rect 76 867 83 873
rect 33 863 47 867
rect 16 856 47 863
rect 16 807 23 856
rect 33 853 47 856
rect 53 833 67 847
rect 73 853 87 867
rect 56 823 63 833
rect 36 816 63 823
rect 36 647 43 816
rect 96 803 103 1073
rect 196 1067 203 1096
rect 213 1093 227 1107
rect 236 1087 243 1133
rect 256 1127 263 1313
rect 296 1303 303 1336
rect 276 1296 303 1303
rect 276 1227 283 1296
rect 316 1287 323 1356
rect 376 1347 383 1433
rect 396 1347 403 1373
rect 416 1347 423 1413
rect 436 1407 443 1553
rect 456 1467 463 1693
rect 476 1607 483 1613
rect 473 1593 487 1607
rect 476 1367 483 1493
rect 373 1333 387 1347
rect 496 1343 503 1633
rect 536 1627 543 1753
rect 656 1747 663 1773
rect 576 1627 583 1633
rect 573 1613 587 1627
rect 513 1603 527 1607
rect 513 1596 543 1603
rect 513 1593 527 1596
rect 536 1563 543 1596
rect 596 1587 603 1633
rect 636 1627 643 1653
rect 636 1587 643 1613
rect 656 1607 663 1713
rect 696 1623 703 1773
rect 716 1647 723 1833
rect 736 1827 743 1993
rect 756 1747 763 2033
rect 776 2007 783 2076
rect 796 2027 803 2093
rect 816 2087 823 2193
rect 836 2087 843 2213
rect 896 2167 903 2273
rect 916 2207 923 2253
rect 936 2227 943 2493
rect 956 2487 963 2513
rect 976 2507 983 2533
rect 1013 2513 1027 2527
rect 1033 2533 1047 2547
rect 1053 2513 1067 2527
rect 956 2307 963 2333
rect 976 2247 983 2433
rect 996 2387 1003 2513
rect 1016 2487 1023 2513
rect 1036 2287 1043 2393
rect 1056 2267 1063 2513
rect 1076 2447 1083 2513
rect 1096 2307 1103 2593
rect 1136 2547 1143 2633
rect 1156 2547 1163 2633
rect 1176 2547 1183 2593
rect 1236 2587 1243 2593
rect 1113 2513 1127 2527
rect 1133 2533 1147 2547
rect 1173 2533 1187 2547
rect 1196 2543 1203 2573
rect 1213 2543 1227 2547
rect 1196 2536 1227 2543
rect 1213 2533 1227 2536
rect 1116 2467 1123 2513
rect 1136 2327 1143 2493
rect 1116 2287 1123 2313
rect 1073 2273 1087 2287
rect 1076 2267 1083 2273
rect 1093 2253 1107 2267
rect 1113 2273 1127 2287
rect 1133 2263 1147 2267
rect 1156 2263 1163 2373
rect 1196 2347 1203 2513
rect 1256 2407 1263 2693
rect 1316 2667 1323 2813
rect 1356 2767 1363 2873
rect 1376 2807 1383 2996
rect 1396 2987 1403 3013
rect 1433 3013 1447 3027
rect 1476 3007 1483 3073
rect 1516 3027 1523 3073
rect 1556 3027 1563 3173
rect 1576 3123 1583 3613
rect 1596 3527 1603 3553
rect 1593 3513 1607 3527
rect 1596 3287 1603 3473
rect 1636 3327 1643 3633
rect 1655 3476 1663 3556
rect 1796 3547 1803 4033
rect 1816 3987 1823 4013
rect 1876 4007 1883 4073
rect 1936 4047 1943 4173
rect 1873 4003 1887 4007
rect 1893 4003 1907 4007
rect 1813 3973 1827 3987
rect 1853 3973 1867 3987
rect 1873 3996 1907 4003
rect 1936 4007 1943 4033
rect 1873 3993 1887 3996
rect 1893 3993 1907 3996
rect 1933 3993 1947 4007
rect 1856 3967 1863 3973
rect 1816 3707 1823 3933
rect 1836 3743 1843 3953
rect 1836 3736 1863 3743
rect 1856 3727 1863 3736
rect 1896 3727 1903 3753
rect 1833 3693 1847 3707
rect 1853 3713 1867 3727
rect 1893 3713 1907 3727
rect 1836 3667 1843 3693
rect 1916 3687 1923 3973
rect 1956 3767 1963 4013
rect 1976 3987 1983 4153
rect 1996 4107 2003 4193
rect 2013 4023 2027 4027
rect 2036 4023 2043 4393
rect 2096 4327 2103 4476
rect 2173 4473 2187 4487
rect 2233 4463 2247 4467
rect 2233 4456 2263 4463
rect 2233 4453 2247 4456
rect 2256 4447 2263 4456
rect 2116 4227 2123 4273
rect 2073 4213 2087 4227
rect 2053 4193 2067 4207
rect 2056 4047 2063 4193
rect 2076 4147 2083 4213
rect 2113 4213 2127 4227
rect 2196 4144 2204 4256
rect 2276 4223 2283 4533
rect 2296 4487 2303 4513
rect 2336 4487 2343 4533
rect 2293 4473 2307 4487
rect 2333 4473 2347 4487
rect 2353 4453 2367 4467
rect 2413 4483 2427 4487
rect 2413 4476 2433 4483
rect 2413 4473 2427 4476
rect 2356 4447 2363 4453
rect 2367 4436 2383 4443
rect 2335 4238 2343 4262
rect 2256 4216 2283 4223
rect 2233 4183 2247 4187
rect 2256 4183 2263 4216
rect 2233 4176 2263 4183
rect 2233 4173 2247 4176
rect 2273 4173 2287 4187
rect 2013 4016 2043 4023
rect 2013 4013 2027 4016
rect 2036 4007 2043 4016
rect 2076 4007 2083 4093
rect 2136 4027 2143 4113
rect 2133 4013 2147 4027
rect 1993 3973 2007 3987
rect 2033 3993 2047 4007
rect 2053 3973 2067 3987
rect 2073 3993 2087 4007
rect 1996 3967 2003 3973
rect 2056 3963 2063 3973
rect 2056 3956 2083 3963
rect 2176 3963 2183 4113
rect 2276 4087 2283 4173
rect 2335 4144 2343 4224
rect 2193 3963 2207 3967
rect 2176 3956 2207 3963
rect 2233 3963 2247 3967
rect 2256 3963 2263 4053
rect 2276 4007 2283 4033
rect 2276 3987 2283 3993
rect 2316 3987 2323 4093
rect 2376 4047 2383 4436
rect 2436 4427 2443 4473
rect 2476 4463 2483 4493
rect 2553 4483 2567 4487
rect 2493 4463 2507 4467
rect 2476 4456 2507 4463
rect 2493 4453 2507 4456
rect 2533 4453 2547 4467
rect 2553 4476 2583 4483
rect 2553 4473 2567 4476
rect 2536 4447 2543 4453
rect 2393 4173 2407 4187
rect 2396 4027 2403 4173
rect 2416 4007 2423 4393
rect 2433 4183 2447 4187
rect 2456 4183 2463 4373
rect 2496 4207 2503 4433
rect 2576 4427 2583 4476
rect 2633 4453 2647 4467
rect 2693 4483 2707 4487
rect 2673 4453 2687 4467
rect 2693 4476 2723 4483
rect 2693 4473 2707 4476
rect 2716 4467 2723 4476
rect 2636 4427 2643 4453
rect 2676 4447 2683 4453
rect 2657 4238 2665 4262
rect 2676 4247 2683 4433
rect 2756 4404 2764 4516
rect 2833 4483 2847 4487
rect 2816 4476 2847 4483
rect 2433 4176 2463 4183
rect 2433 4173 2447 4176
rect 2556 4167 2563 4173
rect 2596 4167 2603 4173
rect 2573 4153 2587 4167
rect 2576 4027 2583 4153
rect 2657 4144 2665 4224
rect 2373 4003 2387 4007
rect 2373 3996 2403 4003
rect 2373 3993 2387 3996
rect 1953 3713 1967 3727
rect 1956 3707 1963 3713
rect 2013 3703 2027 3707
rect 2013 3696 2043 3703
rect 2013 3693 2027 3696
rect 1676 3487 1683 3513
rect 1655 3438 1663 3462
rect 1676 3387 1683 3413
rect 1676 3247 1683 3373
rect 1696 3267 1703 3533
rect 1836 3527 1843 3533
rect 1716 3407 1723 3513
rect 1733 3473 1747 3487
rect 1813 3493 1827 3507
rect 1833 3513 1847 3527
rect 1773 3473 1787 3487
rect 1736 3467 1743 3473
rect 1716 3307 1723 3353
rect 1653 3223 1667 3227
rect 1636 3216 1667 3223
rect 1673 3233 1687 3247
rect 1713 3233 1727 3247
rect 1716 3227 1723 3233
rect 1576 3116 1603 3123
rect 1453 2993 1467 3007
rect 1493 2993 1507 3007
rect 1533 2993 1547 3007
rect 1416 2983 1423 2993
rect 1456 2987 1463 2993
rect 1416 2976 1443 2983
rect 1333 2733 1347 2747
rect 1336 2667 1343 2733
rect 1296 2567 1303 2613
rect 1336 2567 1343 2593
rect 1356 2567 1363 2753
rect 1396 2663 1403 2973
rect 1416 2704 1424 2816
rect 1396 2656 1423 2663
rect 1293 2553 1307 2567
rect 1276 2547 1283 2553
rect 1273 2533 1287 2547
rect 1313 2533 1327 2547
rect 1333 2553 1347 2567
rect 1376 2547 1383 2573
rect 1133 2256 1163 2263
rect 1133 2253 1147 2256
rect 1193 2253 1207 2267
rect 1096 2247 1103 2253
rect 833 2073 847 2087
rect 873 2083 887 2087
rect 896 2083 903 2093
rect 936 2087 943 2113
rect 956 2087 963 2233
rect 1136 2227 1143 2253
rect 853 2053 867 2067
rect 873 2076 903 2083
rect 873 2073 887 2076
rect 896 2067 903 2076
rect 936 2067 943 2073
rect 893 2053 907 2067
rect 933 2053 947 2067
rect 856 2007 863 2053
rect 916 2047 923 2053
rect 953 2033 967 2047
rect 776 1783 783 1913
rect 816 1827 823 1853
rect 836 1807 843 1873
rect 856 1847 863 1953
rect 876 1867 883 2033
rect 896 1987 903 2013
rect 896 1807 903 1873
rect 936 1863 943 2013
rect 956 1887 963 2033
rect 976 2007 983 2213
rect 996 2067 1003 2073
rect 1016 2067 1023 2093
rect 1036 2067 1043 2113
rect 1116 2087 1123 2093
rect 1156 2087 1163 2213
rect 993 2053 1007 2067
rect 1033 2053 1047 2067
rect 1053 2043 1067 2047
rect 1076 2043 1083 2073
rect 1053 2036 1083 2043
rect 1116 2047 1123 2073
rect 1053 2033 1067 2036
rect 1113 2033 1127 2047
rect 996 1987 1003 2013
rect 916 1856 943 1863
rect 916 1827 923 1856
rect 776 1776 803 1783
rect 676 1616 703 1623
rect 553 1573 567 1587
rect 593 1573 607 1587
rect 633 1573 647 1587
rect 393 1293 407 1307
rect 453 1323 467 1327
rect 476 1336 503 1343
rect 516 1556 543 1563
rect 476 1323 483 1336
rect 516 1327 523 1556
rect 536 1327 543 1533
rect 556 1527 563 1573
rect 453 1316 483 1323
rect 453 1313 467 1316
rect 433 1293 447 1307
rect 296 1207 303 1273
rect 336 1187 343 1293
rect 296 1147 303 1173
rect 356 1147 363 1273
rect 376 1187 383 1293
rect 396 1167 403 1293
rect 436 1247 443 1293
rect 456 1227 463 1313
rect 476 1167 483 1293
rect 553 1293 567 1307
rect 556 1287 563 1293
rect 513 1273 527 1287
rect 376 1143 383 1153
rect 376 1136 403 1143
rect 296 1103 303 1113
rect 313 1103 327 1107
rect 233 1073 247 1087
rect 296 1096 327 1103
rect 313 1093 327 1096
rect 353 1093 367 1107
rect 133 863 147 867
rect 176 863 183 1053
rect 256 867 263 1053
rect 296 887 303 1073
rect 356 1067 363 1093
rect 396 1087 403 1136
rect 416 1127 423 1153
rect 416 1107 423 1113
rect 436 1107 443 1133
rect 413 1093 427 1107
rect 436 1087 443 1093
rect 433 1073 447 1087
rect 496 1067 503 1273
rect 516 1227 523 1273
rect 576 1247 583 1573
rect 616 1567 623 1573
rect 653 1553 667 1567
rect 656 1547 663 1553
rect 593 1293 607 1307
rect 633 1293 647 1307
rect 596 1287 603 1293
rect 596 1267 603 1273
rect 556 1147 563 1193
rect 576 1127 583 1213
rect 616 1207 623 1273
rect 636 1247 643 1293
rect 656 1187 663 1313
rect 573 1113 587 1127
rect 527 1076 533 1083
rect 133 856 163 863
rect 176 856 203 863
rect 133 853 147 856
rect 96 796 123 803
rect 33 643 47 647
rect 16 636 47 643
rect 116 647 123 796
rect 136 667 143 813
rect 156 807 163 856
rect 196 827 203 856
rect 213 833 227 847
rect 173 813 187 827
rect 176 787 183 813
rect 216 707 223 833
rect 273 813 287 827
rect 296 823 303 873
rect 376 847 383 853
rect 313 823 327 827
rect 296 816 327 823
rect 156 667 163 673
rect 153 653 167 667
rect 73 643 87 647
rect 16 387 23 636
rect 33 633 47 636
rect 73 636 103 643
rect 73 633 87 636
rect 96 407 103 636
rect 113 633 127 647
rect 173 613 187 627
rect 213 613 227 627
rect 96 387 103 393
rect 156 387 163 613
rect 176 607 183 613
rect 196 403 203 613
rect 216 607 223 613
rect 236 427 243 633
rect 176 396 203 403
rect 13 373 27 387
rect 53 383 67 387
rect 33 353 47 367
rect 53 376 83 383
rect 53 373 67 376
rect 36 207 43 353
rect 76 327 83 376
rect 93 373 107 387
rect 133 383 147 387
rect 113 353 127 367
rect 133 376 153 383
rect 133 373 147 376
rect 36 163 43 193
rect 36 156 63 163
rect 56 147 63 156
rect 76 147 83 173
rect 96 167 103 333
rect 116 187 123 353
rect 176 347 183 396
rect 236 387 243 393
rect 233 373 247 387
rect 256 367 263 693
rect 276 667 283 813
rect 296 787 303 816
rect 313 813 327 816
rect 373 833 387 847
rect 396 723 403 813
rect 376 716 403 723
rect 316 667 323 673
rect 313 653 327 667
rect 356 647 363 673
rect 376 667 383 716
rect 416 707 423 873
rect 433 813 447 827
rect 436 807 443 813
rect 356 627 363 633
rect 396 627 403 693
rect 293 613 307 627
rect 353 613 367 627
rect 296 607 303 613
rect 276 387 283 573
rect 316 527 323 613
rect 413 593 427 607
rect 316 387 323 453
rect 273 373 287 387
rect 293 353 307 367
rect 313 373 327 387
rect 296 347 303 353
rect 256 327 263 333
rect 136 187 143 193
rect 133 173 147 187
rect 96 147 103 153
rect 53 133 67 147
rect 93 133 107 147
rect 236 147 243 193
rect 316 187 323 333
rect 336 187 343 413
rect 356 387 363 493
rect 396 367 403 433
rect 416 407 423 593
rect 436 507 443 673
rect 456 667 463 853
rect 496 847 503 893
rect 516 847 523 913
rect 513 833 527 847
rect 473 813 487 827
rect 476 747 483 813
rect 536 747 543 1053
rect 556 763 563 1033
rect 576 907 583 1073
rect 576 847 583 853
rect 596 847 603 1173
rect 573 833 587 847
rect 616 823 623 1173
rect 656 1107 663 1153
rect 676 1123 683 1616
rect 756 1607 763 1693
rect 733 1573 747 1587
rect 753 1593 767 1607
rect 696 1507 703 1553
rect 716 1387 723 1573
rect 736 1527 743 1573
rect 736 1347 743 1453
rect 693 1293 707 1307
rect 753 1313 767 1327
rect 696 1267 703 1293
rect 756 1287 763 1313
rect 716 1227 723 1273
rect 716 1127 723 1193
rect 736 1127 743 1173
rect 776 1143 783 1633
rect 796 1607 803 1776
rect 833 1793 847 1807
rect 893 1793 907 1807
rect 933 1793 947 1807
rect 936 1787 943 1793
rect 913 1773 927 1787
rect 816 1727 823 1753
rect 856 1727 863 1753
rect 816 1587 823 1613
rect 876 1607 883 1753
rect 916 1747 923 1773
rect 936 1707 943 1773
rect 956 1747 963 1853
rect 1016 1847 1023 1893
rect 1036 1867 1043 2013
rect 1036 1847 1043 1853
rect 1056 1827 1063 2013
rect 1013 1793 1027 1807
rect 1076 1803 1083 1993
rect 1096 1847 1103 2013
rect 1176 2007 1183 2253
rect 1196 2247 1203 2253
rect 1256 2227 1263 2293
rect 1233 2053 1247 2067
rect 1276 2067 1283 2493
rect 1316 2347 1323 2533
rect 1353 2513 1367 2527
rect 1373 2533 1387 2547
rect 1393 2513 1407 2527
rect 1356 2487 1363 2513
rect 1396 2507 1403 2513
rect 1416 2507 1423 2656
rect 1436 2587 1443 2976
rect 1496 2927 1503 2993
rect 1536 2987 1543 2993
rect 1456 2767 1463 2913
rect 1556 2867 1563 2993
rect 1456 2587 1463 2753
rect 1493 2733 1507 2747
rect 1533 2743 1547 2747
rect 1556 2743 1563 2853
rect 1576 2847 1583 2973
rect 1596 2967 1603 3116
rect 1616 3047 1623 3153
rect 1533 2736 1563 2743
rect 1533 2733 1547 2736
rect 1456 2567 1463 2573
rect 1476 2567 1483 2673
rect 1496 2607 1503 2733
rect 1453 2553 1467 2567
rect 1496 2543 1503 2573
rect 1476 2536 1503 2543
rect 1296 2224 1304 2336
rect 1316 2183 1323 2313
rect 1333 2253 1347 2267
rect 1336 2247 1343 2253
rect 1296 2176 1323 2183
rect 1296 2107 1303 2176
rect 1316 2107 1323 2133
rect 1313 2093 1327 2107
rect 1096 1807 1103 1813
rect 1056 1796 1083 1803
rect 1016 1787 1023 1793
rect 1036 1747 1043 1773
rect 916 1627 923 1633
rect 956 1607 963 1613
rect 893 1573 907 1587
rect 953 1593 967 1607
rect 876 1543 883 1573
rect 896 1567 903 1573
rect 856 1536 883 1543
rect 796 1347 803 1493
rect 796 1227 803 1293
rect 816 1287 823 1413
rect 836 1367 843 1473
rect 856 1467 863 1536
rect 896 1527 903 1553
rect 916 1507 923 1573
rect 853 1293 867 1307
rect 756 1136 783 1143
rect 676 1116 703 1123
rect 633 1073 647 1087
rect 653 1093 667 1107
rect 636 1027 643 1073
rect 696 887 703 1116
rect 713 1113 727 1127
rect 756 927 763 1136
rect 776 1027 783 1073
rect 776 867 783 993
rect 656 847 663 853
rect 696 847 703 853
rect 633 823 647 827
rect 616 816 647 823
rect 653 833 667 847
rect 713 843 727 847
rect 713 836 743 843
rect 713 833 727 836
rect 633 813 647 816
rect 593 793 607 807
rect 596 767 603 793
rect 556 756 583 763
rect 436 407 443 473
rect 456 407 463 653
rect 536 647 543 713
rect 513 613 527 627
rect 533 633 547 647
rect 516 603 523 613
rect 516 596 543 603
rect 476 403 483 513
rect 496 487 503 593
rect 536 587 543 596
rect 516 507 523 573
rect 556 567 563 733
rect 576 663 583 756
rect 616 667 623 693
rect 576 656 603 663
rect 476 396 503 403
rect 353 333 367 347
rect 356 327 363 333
rect 436 327 443 393
rect 456 387 463 393
rect 496 387 503 396
rect 473 353 487 367
rect 476 327 483 353
rect 516 327 523 453
rect 596 427 603 656
rect 616 647 623 653
rect 636 647 643 793
rect 613 633 627 647
rect 656 627 663 753
rect 676 687 683 793
rect 696 663 703 773
rect 676 656 703 663
rect 676 647 683 656
rect 716 647 723 793
rect 736 767 743 836
rect 753 833 767 847
rect 773 853 787 867
rect 756 827 763 833
rect 673 633 687 647
rect 653 613 667 627
rect 693 613 707 627
rect 536 387 543 413
rect 533 373 547 387
rect 573 373 587 387
rect 553 353 567 367
rect 356 287 363 313
rect 476 307 483 313
rect 256 167 263 173
rect 356 167 363 253
rect 253 153 267 167
rect 233 133 247 147
rect 353 153 367 167
rect 376 147 383 153
rect 373 133 387 147
rect 76 127 83 133
rect 73 113 87 127
rect 416 123 423 233
rect 436 187 443 293
rect 556 267 563 353
rect 576 343 583 373
rect 576 336 603 343
rect 433 123 447 127
rect 416 116 447 123
rect 476 127 483 173
rect 496 147 503 153
rect 493 133 507 147
rect 433 113 447 116
rect 473 113 487 127
rect 536 127 543 173
rect 556 147 563 193
rect 596 187 603 336
rect 616 207 623 493
rect 636 447 643 613
rect 696 547 703 613
rect 656 367 663 393
rect 696 367 703 393
rect 633 333 647 347
rect 653 353 667 367
rect 673 333 687 347
rect 693 353 707 367
rect 636 327 643 333
rect 676 227 683 333
rect 696 203 703 313
rect 736 247 743 753
rect 776 663 783 733
rect 796 687 803 1193
rect 816 1127 823 1273
rect 836 1167 843 1293
rect 856 1287 863 1293
rect 876 1263 883 1453
rect 936 1427 943 1573
rect 856 1256 883 1263
rect 856 1247 863 1256
rect 836 1107 843 1133
rect 856 1127 863 1213
rect 876 1107 883 1233
rect 896 1227 903 1353
rect 956 1347 963 1373
rect 976 1367 983 1673
rect 996 1587 1003 1633
rect 1016 1607 1023 1733
rect 1056 1603 1063 1796
rect 1093 1793 1107 1807
rect 1116 1763 1123 1993
rect 1147 1856 1153 1863
rect 1196 1827 1203 2053
rect 1133 1803 1147 1807
rect 1133 1796 1163 1803
rect 1133 1793 1147 1796
rect 1156 1787 1163 1796
rect 1173 1793 1187 1807
rect 1193 1813 1207 1827
rect 1096 1756 1123 1763
rect 1076 1627 1083 1753
rect 1056 1596 1083 1603
rect 993 1573 1007 1587
rect 1033 1583 1047 1587
rect 1027 1576 1047 1583
rect 1033 1573 1047 1576
rect 1076 1543 1083 1596
rect 1096 1567 1103 1756
rect 1136 1667 1143 1773
rect 1176 1747 1183 1793
rect 1116 1587 1123 1633
rect 1136 1607 1143 1653
rect 1133 1593 1147 1607
rect 1196 1587 1203 1593
rect 1216 1587 1223 2053
rect 1236 1847 1243 2053
rect 1276 1847 1283 2033
rect 1296 1847 1303 2013
rect 1233 1793 1247 1807
rect 1236 1767 1243 1793
rect 1256 1727 1263 1813
rect 1273 1793 1287 1807
rect 1276 1747 1283 1793
rect 1256 1647 1263 1673
rect 1193 1573 1207 1587
rect 1276 1567 1283 1693
rect 1296 1687 1303 1773
rect 1316 1707 1323 2053
rect 1356 2043 1363 2333
rect 1416 2267 1423 2473
rect 1436 2427 1443 2533
rect 1476 2367 1483 2536
rect 1435 2318 1443 2342
rect 1373 2253 1387 2267
rect 1376 2207 1383 2253
rect 1416 2107 1423 2253
rect 1435 2224 1443 2304
rect 1476 2223 1483 2333
rect 1496 2283 1503 2373
rect 1576 2347 1583 2833
rect 1616 2827 1623 2953
rect 1596 2704 1604 2816
rect 1636 2787 1643 3216
rect 1653 3213 1667 3216
rect 1716 3207 1723 3213
rect 1656 3047 1663 3093
rect 1696 3047 1703 3153
rect 1736 3147 1743 3353
rect 1653 3033 1667 3047
rect 1673 3013 1687 3027
rect 1693 3033 1707 3047
rect 1716 3027 1723 3073
rect 1713 3013 1727 3027
rect 1633 2733 1647 2747
rect 1636 2707 1643 2733
rect 1656 2667 1663 2973
rect 1676 2887 1683 3013
rect 1696 2927 1703 2993
rect 1736 2983 1743 3113
rect 1756 3107 1763 3453
rect 1776 3407 1783 3473
rect 1816 3467 1823 3493
rect 1796 3303 1803 3373
rect 1787 3296 1803 3303
rect 1816 3247 1823 3273
rect 1836 3267 1843 3293
rect 1856 3267 1863 3433
rect 1876 3423 1883 3673
rect 1916 3527 1923 3633
rect 1893 3493 1907 3507
rect 1913 3513 1927 3527
rect 1896 3487 1903 3493
rect 1896 3447 1903 3473
rect 1876 3416 1903 3423
rect 1896 3287 1903 3416
rect 1853 3253 1867 3267
rect 1773 3233 1787 3247
rect 1776 3167 1783 3233
rect 1813 3233 1827 3247
rect 1873 3233 1887 3247
rect 1876 3227 1883 3233
rect 1876 3207 1883 3213
rect 1796 3047 1803 3153
rect 1816 3047 1823 3133
rect 1793 3033 1807 3047
rect 1836 3007 1843 3193
rect 1896 3123 1903 3213
rect 1916 3147 1923 3473
rect 1936 3367 1943 3613
rect 1956 3487 1963 3673
rect 1996 3507 2003 3593
rect 2036 3523 2043 3696
rect 2076 3683 2083 3956
rect 2193 3953 2207 3956
rect 2233 3956 2263 3963
rect 2273 3973 2287 3987
rect 2313 3973 2327 3987
rect 2296 3967 2303 3973
rect 2233 3953 2247 3956
rect 2293 3953 2307 3967
rect 2333 3953 2347 3967
rect 2336 3763 2343 3953
rect 2316 3756 2343 3763
rect 2093 3703 2107 3707
rect 2093 3696 2123 3703
rect 2093 3693 2107 3696
rect 2076 3676 2103 3683
rect 2053 3523 2067 3527
rect 2036 3516 2067 3523
rect 2013 3483 2027 3487
rect 2036 3483 2043 3516
rect 2053 3513 2067 3516
rect 2013 3476 2043 3483
rect 2013 3473 2027 3476
rect 2073 3473 2087 3487
rect 1956 3247 1963 3273
rect 1976 3267 1983 3373
rect 1953 3233 1967 3247
rect 1993 3233 2007 3247
rect 1973 3213 1987 3227
rect 1896 3116 1923 3123
rect 1856 3047 1863 3093
rect 1876 3067 1883 3093
rect 1873 3053 1887 3067
rect 1853 3033 1867 3047
rect 1716 2976 1743 2983
rect 1696 2827 1703 2893
rect 1673 2743 1687 2747
rect 1696 2743 1703 2813
rect 1673 2736 1703 2743
rect 1673 2733 1687 2736
rect 1696 2687 1703 2736
rect 1596 2527 1603 2593
rect 1513 2283 1527 2287
rect 1496 2276 1527 2283
rect 1513 2273 1527 2276
rect 1533 2253 1547 2267
rect 1536 2227 1543 2253
rect 1576 2247 1583 2253
rect 1456 2216 1483 2223
rect 1436 2083 1443 2093
rect 1416 2076 1443 2083
rect 1376 2067 1383 2073
rect 1416 2067 1423 2076
rect 1356 2036 1383 2043
rect 1356 1987 1363 2013
rect 1353 1803 1367 1807
rect 1376 1803 1383 2036
rect 1393 2033 1407 2047
rect 1413 2053 1427 2067
rect 1396 2027 1403 2033
rect 1456 1927 1463 2216
rect 1556 2067 1563 2073
rect 1473 2033 1487 2047
rect 1513 2033 1527 2047
rect 1553 2053 1567 2067
rect 1573 2033 1587 2047
rect 1476 2027 1483 2033
rect 1516 2007 1523 2033
rect 1576 2007 1583 2033
rect 1336 1796 1383 1803
rect 1336 1627 1343 1796
rect 1353 1793 1367 1796
rect 1373 1753 1387 1767
rect 1376 1727 1383 1753
rect 1356 1607 1363 1653
rect 1293 1583 1307 1587
rect 1293 1576 1323 1583
rect 1293 1573 1307 1576
rect 1253 1553 1267 1567
rect 1056 1536 1083 1543
rect 996 1507 1003 1533
rect 1036 1447 1043 1533
rect 953 1333 967 1347
rect 993 1313 1007 1327
rect 916 1287 923 1293
rect 996 1287 1003 1313
rect 813 1073 827 1087
rect 833 1093 847 1107
rect 873 1093 887 1107
rect 856 1087 863 1093
rect 853 1073 867 1087
rect 816 1027 823 1073
rect 896 1067 903 1153
rect 916 1107 923 1273
rect 996 1207 1003 1253
rect 976 1127 983 1153
rect 996 1127 1003 1193
rect 1036 1187 1043 1333
rect 1056 1267 1063 1536
rect 1096 1367 1103 1533
rect 1133 1313 1147 1327
rect 1036 1127 1043 1133
rect 913 1093 927 1107
rect 953 1093 967 1107
rect 973 1113 987 1127
rect 993 1113 1007 1127
rect 1013 1093 1027 1107
rect 1033 1113 1047 1127
rect 1056 1123 1063 1193
rect 1096 1167 1103 1293
rect 1056 1116 1083 1123
rect 956 1087 963 1093
rect 816 707 823 913
rect 836 867 843 973
rect 856 867 863 893
rect 853 853 867 867
rect 776 656 803 663
rect 796 647 803 656
rect 753 643 767 647
rect 753 636 783 643
rect 753 633 767 636
rect 776 607 783 636
rect 793 633 807 647
rect 776 367 783 533
rect 836 403 843 653
rect 856 647 863 813
rect 876 787 883 1053
rect 896 987 903 1033
rect 896 867 903 933
rect 916 867 923 893
rect 913 853 927 867
rect 933 833 947 847
rect 936 807 943 833
rect 976 827 983 853
rect 996 727 1003 953
rect 1016 927 1023 1093
rect 1076 967 1083 1116
rect 1076 887 1083 933
rect 1096 867 1103 1153
rect 1116 1147 1123 1313
rect 1136 1207 1143 1313
rect 1156 1307 1163 1553
rect 1176 1447 1183 1553
rect 1256 1547 1263 1553
rect 1196 1487 1203 1533
rect 1236 1507 1243 1533
rect 1296 1527 1303 1553
rect 1316 1507 1323 1576
rect 1353 1593 1367 1607
rect 1176 1327 1183 1333
rect 1196 1327 1203 1373
rect 1173 1313 1187 1327
rect 1193 1273 1207 1287
rect 1196 1247 1203 1273
rect 1196 1227 1203 1233
rect 1216 1187 1223 1353
rect 1256 1347 1263 1393
rect 1253 1333 1267 1347
rect 1233 1293 1247 1307
rect 1136 1127 1143 1153
rect 1176 1127 1183 1173
rect 1133 1113 1147 1127
rect 1116 1107 1123 1113
rect 1113 1093 1127 1107
rect 1153 1093 1167 1107
rect 1173 1113 1187 1127
rect 1156 1087 1163 1093
rect 1156 987 1163 1073
rect 1116 867 1123 913
rect 1116 847 1123 853
rect 1033 833 1047 847
rect 1073 833 1087 847
rect 1036 767 1043 833
rect 876 647 883 653
rect 873 633 887 647
rect 896 627 903 693
rect 916 647 923 673
rect 956 647 963 693
rect 913 633 927 647
rect 953 633 967 647
rect 856 407 863 593
rect 876 467 883 593
rect 896 587 903 613
rect 876 443 883 453
rect 876 436 903 443
rect 816 396 843 403
rect 753 333 767 347
rect 816 347 823 396
rect 876 387 883 413
rect 896 387 903 436
rect 936 387 943 393
rect 853 353 867 367
rect 873 373 887 387
rect 913 353 927 367
rect 933 373 947 387
rect 756 307 763 333
rect 793 333 807 347
rect 796 327 803 333
rect 773 313 787 327
rect 776 203 783 313
rect 816 227 823 293
rect 856 227 863 353
rect 916 327 923 353
rect 916 267 923 313
rect 956 287 963 353
rect 896 227 903 233
rect 676 196 703 203
rect 756 196 803 203
rect 533 113 547 127
rect 596 127 603 153
rect 676 167 683 196
rect 756 187 763 196
rect 796 187 803 196
rect 816 187 823 213
rect 813 173 827 187
rect 613 133 627 147
rect 653 133 667 147
rect 673 153 687 167
rect 573 113 587 127
rect 576 103 583 113
rect 616 107 623 133
rect 656 127 663 133
rect 836 107 843 133
rect 576 96 593 103
rect 856 47 863 193
rect 876 127 883 153
rect 896 147 903 213
rect 976 207 983 433
rect 996 427 1003 653
rect 1016 647 1023 673
rect 1056 667 1063 833
rect 1076 787 1083 833
rect 1113 833 1127 847
rect 1153 843 1167 847
rect 1176 843 1183 953
rect 1196 947 1203 1153
rect 1236 1147 1243 1293
rect 1256 1267 1263 1293
rect 1253 1073 1267 1087
rect 1256 967 1263 1073
rect 1196 847 1203 913
rect 1216 887 1223 893
rect 1276 887 1283 1333
rect 1336 1327 1343 1553
rect 1376 1367 1383 1613
rect 1396 1407 1403 1913
rect 1436 1827 1443 1873
rect 1576 1827 1583 1993
rect 1436 1807 1443 1813
rect 1433 1793 1447 1807
rect 1453 1773 1467 1787
rect 1513 1793 1527 1807
rect 1573 1813 1587 1827
rect 1516 1787 1523 1793
rect 1493 1773 1507 1787
rect 1456 1747 1463 1773
rect 1496 1767 1503 1773
rect 1536 1647 1543 1793
rect 1433 1623 1447 1627
rect 1433 1616 1463 1623
rect 1433 1613 1447 1616
rect 1456 1587 1463 1616
rect 1453 1583 1467 1587
rect 1436 1576 1467 1583
rect 1416 1487 1423 1553
rect 1436 1507 1443 1576
rect 1453 1573 1467 1576
rect 1476 1567 1483 1633
rect 1576 1627 1583 1633
rect 1596 1627 1603 2493
rect 1616 2484 1624 2596
rect 1656 2567 1663 2613
rect 1653 2553 1667 2567
rect 1636 2387 1643 2533
rect 1616 1827 1623 2273
rect 1636 2224 1644 2336
rect 1656 2267 1663 2513
rect 1676 2487 1683 2633
rect 1696 2567 1703 2673
rect 1716 2483 1723 2976
rect 1796 2947 1803 2993
rect 1735 2798 1743 2822
rect 1756 2807 1763 2873
rect 1735 2704 1743 2784
rect 1776 2687 1783 2793
rect 1836 2787 1843 2973
rect 1793 2733 1807 2747
rect 1796 2607 1803 2733
rect 1856 2707 1863 2733
rect 1696 2476 1723 2483
rect 1673 2253 1687 2267
rect 1676 2227 1683 2253
rect 1696 2187 1703 2476
rect 1713 2263 1727 2267
rect 1736 2263 1743 2553
rect 1755 2516 1763 2596
rect 1773 2553 1787 2567
rect 1755 2478 1763 2502
rect 1776 2427 1783 2553
rect 1836 2547 1843 2653
rect 1833 2533 1847 2547
rect 1853 2513 1867 2527
rect 1816 2507 1823 2513
rect 1856 2487 1863 2513
rect 1876 2483 1883 3013
rect 1916 2847 1923 3116
rect 1936 3067 1943 3193
rect 1976 3147 1983 3213
rect 1996 3187 2003 3233
rect 2016 3163 2023 3453
rect 2036 3243 2043 3273
rect 2076 3267 2083 3473
rect 2096 3467 2103 3676
rect 2116 3547 2123 3696
rect 2156 3607 2163 3733
rect 2316 3727 2323 3756
rect 2336 3727 2343 3733
rect 2193 3723 2207 3727
rect 2176 3716 2207 3723
rect 2176 3587 2183 3716
rect 2193 3713 2207 3716
rect 2333 3713 2347 3727
rect 2176 3567 2183 3573
rect 2156 3507 2163 3513
rect 2133 3473 2147 3487
rect 2153 3493 2167 3507
rect 2213 3503 2227 3507
rect 2173 3483 2187 3487
rect 2196 3496 2227 3503
rect 2196 3483 2203 3496
rect 2173 3476 2203 3483
rect 2213 3493 2227 3496
rect 2236 3487 2243 3513
rect 2173 3473 2187 3476
rect 2233 3473 2247 3487
rect 2273 3473 2287 3487
rect 2096 3247 2103 3413
rect 2116 3267 2123 3473
rect 2136 3463 2143 3473
rect 2136 3456 2163 3463
rect 2156 3347 2163 3456
rect 2136 3247 2143 3313
rect 2156 3247 2163 3333
rect 2053 3243 2067 3247
rect 2036 3236 2067 3243
rect 2053 3233 2067 3236
rect 2093 3233 2107 3247
rect 1996 3156 2023 3163
rect 1956 3067 1963 3113
rect 1953 3053 1967 3067
rect 1996 3047 2003 3156
rect 2036 3143 2043 3213
rect 2016 3136 2043 3143
rect 1933 3013 1947 3027
rect 1973 3013 1987 3027
rect 1993 3033 2007 3047
rect 1896 2767 1903 2793
rect 1936 2787 1943 3013
rect 1976 3007 1983 3013
rect 2016 2967 2023 3136
rect 2036 3067 2043 3093
rect 2033 3053 2047 3067
rect 2076 3027 2083 3193
rect 2096 3047 2103 3073
rect 2116 3067 2123 3213
rect 2133 3193 2147 3207
rect 2136 3087 2143 3193
rect 2093 3033 2107 3047
rect 2156 3027 2163 3113
rect 2176 3107 2183 3473
rect 2276 3307 2283 3473
rect 2276 3227 2283 3273
rect 2296 3267 2303 3553
rect 2316 3547 2323 3593
rect 2313 3533 2327 3547
rect 2356 3367 2363 3993
rect 2376 3707 2383 3913
rect 2396 3683 2403 3996
rect 2413 3993 2427 4007
rect 2376 3676 2403 3683
rect 2376 3627 2383 3676
rect 2416 3664 2424 3776
rect 2396 3543 2403 3653
rect 2436 3567 2443 4013
rect 2473 3973 2487 3987
rect 2476 3907 2483 3973
rect 2476 3747 2483 3893
rect 2555 3758 2563 3782
rect 2453 3693 2467 3707
rect 2456 3687 2463 3693
rect 2396 3536 2423 3543
rect 2336 3247 2343 3293
rect 2356 3267 2363 3273
rect 2396 3267 2403 3293
rect 2353 3253 2367 3267
rect 2313 3243 2327 3247
rect 2296 3236 2327 3243
rect 2213 3063 2227 3067
rect 2213 3056 2263 3063
rect 2213 3053 2227 3056
rect 1976 2767 1983 2773
rect 2016 2767 2023 2793
rect 1913 2763 1927 2767
rect 1913 2756 1933 2763
rect 1913 2753 1927 2756
rect 1936 2743 1943 2753
rect 1953 2743 1967 2747
rect 1936 2736 1967 2743
rect 1973 2753 1987 2767
rect 1953 2733 1967 2736
rect 2013 2753 2027 2767
rect 2033 2733 2047 2747
rect 1916 2547 1923 2673
rect 1936 2567 1943 2713
rect 1893 2513 1907 2527
rect 1913 2533 1927 2547
rect 1933 2513 1947 2527
rect 1896 2507 1903 2513
rect 1876 2476 1903 2483
rect 1775 2318 1783 2342
rect 1713 2256 1743 2263
rect 1713 2253 1727 2256
rect 1716 2207 1723 2253
rect 1775 2224 1783 2304
rect 1796 2267 1803 2473
rect 1816 2207 1823 2453
rect 1853 2283 1867 2287
rect 1836 2276 1867 2283
rect 1836 2247 1843 2276
rect 1853 2273 1867 2276
rect 1873 2233 1887 2247
rect 1876 2227 1883 2233
rect 1636 2067 1643 2173
rect 1656 2087 1663 2113
rect 1696 2087 1703 2153
rect 1756 2107 1763 2133
rect 1653 2073 1667 2087
rect 1776 2087 1783 2173
rect 1816 2087 1823 2153
rect 1836 2107 1843 2153
rect 1833 2093 1847 2107
rect 1773 2073 1787 2087
rect 1813 2073 1827 2087
rect 1856 2087 1863 2093
rect 1853 2073 1867 2087
rect 1613 1753 1627 1767
rect 1616 1687 1623 1753
rect 1573 1613 1587 1627
rect 1473 1553 1487 1567
rect 1313 1293 1327 1307
rect 1373 1313 1387 1327
rect 1353 1293 1367 1307
rect 1296 1147 1303 1293
rect 1316 1287 1323 1293
rect 1313 1073 1327 1087
rect 1316 1067 1323 1073
rect 1216 867 1223 873
rect 1213 853 1227 867
rect 1153 836 1183 843
rect 1153 833 1167 836
rect 1253 853 1267 867
rect 1256 847 1263 853
rect 1296 847 1303 1013
rect 1316 847 1323 913
rect 1336 867 1343 1253
rect 1356 1207 1363 1293
rect 1376 1267 1383 1313
rect 1396 1243 1403 1353
rect 1376 1236 1403 1243
rect 1356 1127 1363 1133
rect 1376 1127 1383 1236
rect 1353 1113 1367 1127
rect 1396 1107 1403 1213
rect 1416 1127 1423 1393
rect 1436 1387 1443 1413
rect 1456 1347 1463 1493
rect 1476 1327 1483 1373
rect 1496 1367 1503 1473
rect 1516 1347 1523 1433
rect 1536 1427 1543 1613
rect 1593 1573 1607 1587
rect 1636 1583 1643 1753
rect 1656 1747 1663 1973
rect 1716 1907 1723 2053
rect 1736 2027 1743 2053
rect 1876 2007 1883 2153
rect 1896 2127 1903 2476
rect 1936 2427 1943 2513
rect 1956 2487 1963 2693
rect 2036 2687 2043 2733
rect 2056 2707 2063 2793
rect 2076 2647 2083 2993
rect 2216 2787 2223 3013
rect 2256 2847 2263 3056
rect 2093 2733 2107 2747
rect 2096 2727 2103 2733
rect 2156 2743 2163 2753
rect 2173 2743 2187 2747
rect 2156 2736 2187 2743
rect 2213 2743 2227 2747
rect 2236 2743 2243 2793
rect 2276 2767 2283 3073
rect 2296 3047 2303 3236
rect 2313 3233 2327 3236
rect 2373 3233 2387 3247
rect 2393 3253 2407 3267
rect 2376 3147 2383 3233
rect 2356 3047 2363 3093
rect 2396 3047 2403 3213
rect 2393 3033 2407 3047
rect 2416 3043 2423 3536
rect 2436 3523 2443 3533
rect 2453 3523 2467 3527
rect 2436 3516 2467 3523
rect 2436 3067 2443 3516
rect 2453 3513 2467 3516
rect 2477 3476 2485 3556
rect 2477 3438 2485 3462
rect 2477 3278 2485 3302
rect 2477 3184 2485 3264
rect 2456 3087 2463 3173
rect 2456 3067 2463 3073
rect 2453 3053 2467 3067
rect 2416 3036 2443 3043
rect 2396 2983 2403 2993
rect 2396 2976 2423 2983
rect 2173 2733 2187 2736
rect 2113 2713 2127 2727
rect 2213 2736 2243 2743
rect 2213 2733 2227 2736
rect 2253 2733 2267 2747
rect 2256 2727 2263 2733
rect 2293 2733 2307 2747
rect 2273 2713 2287 2727
rect 2116 2687 2123 2713
rect 2276 2707 2283 2713
rect 2296 2687 2303 2733
rect 2096 2587 2103 2673
rect 2196 2587 2203 2633
rect 2093 2573 2107 2587
rect 2193 2573 2207 2587
rect 1976 2547 1983 2573
rect 2076 2567 2083 2573
rect 2073 2553 2087 2567
rect 1973 2533 1987 2547
rect 2033 2513 2047 2527
rect 2036 2507 2043 2513
rect 1976 2287 1983 2293
rect 1953 2253 1967 2267
rect 1993 2263 2007 2267
rect 2036 2263 2043 2473
rect 1993 2256 2043 2263
rect 1993 2253 2007 2256
rect 1933 2233 1947 2247
rect 1956 2243 1963 2253
rect 1956 2236 1983 2243
rect 1916 2127 1923 2233
rect 1936 2207 1943 2233
rect 1936 2167 1943 2193
rect 1916 2087 1923 2113
rect 1956 2107 1963 2213
rect 1976 2127 1983 2236
rect 1936 2087 1943 2093
rect 1976 2087 1983 2113
rect 1996 2087 2003 2173
rect 2056 2147 2063 2513
rect 2096 2467 2103 2533
rect 2136 2523 2143 2573
rect 2233 2563 2247 2567
rect 2216 2556 2247 2563
rect 2276 2567 2283 2653
rect 2216 2547 2223 2556
rect 2233 2553 2247 2556
rect 2273 2553 2287 2567
rect 2116 2516 2143 2523
rect 1933 2073 1947 2087
rect 1913 2063 1927 2067
rect 1896 2056 1927 2063
rect 1896 2027 1903 2056
rect 1913 2053 1927 2056
rect 1973 2073 1987 2087
rect 1993 2073 2007 2087
rect 2013 2053 2027 2067
rect 2056 2067 2063 2113
rect 2076 2083 2083 2293
rect 2096 2224 2104 2336
rect 2116 2227 2123 2516
rect 2133 2253 2147 2267
rect 2136 2087 2143 2253
rect 2156 2147 2163 2413
rect 2173 2253 2187 2267
rect 2176 2203 2183 2253
rect 2196 2227 2203 2533
rect 2235 2318 2243 2342
rect 2176 2196 2203 2203
rect 2176 2087 2183 2173
rect 2076 2076 2103 2083
rect 2096 2067 2103 2076
rect 2133 2073 2147 2087
rect 2116 2067 2123 2073
rect 2053 2063 2067 2067
rect 2053 2056 2083 2063
rect 2053 2053 2067 2056
rect 1896 1983 1903 2013
rect 1876 1976 1903 1983
rect 1676 1627 1683 1813
rect 1716 1807 1723 1833
rect 1756 1827 1763 1893
rect 1876 1827 1883 1976
rect 1753 1813 1767 1827
rect 1693 1773 1707 1787
rect 1873 1823 1887 1827
rect 1773 1793 1787 1807
rect 1813 1793 1827 1807
rect 1856 1816 1887 1823
rect 1696 1707 1703 1773
rect 1653 1583 1667 1587
rect 1636 1576 1667 1583
rect 1556 1467 1563 1573
rect 1556 1347 1563 1393
rect 1473 1313 1487 1327
rect 1553 1333 1567 1347
rect 1493 1293 1507 1307
rect 1436 1223 1443 1293
rect 1496 1287 1503 1293
rect 1536 1267 1543 1313
rect 1436 1216 1463 1223
rect 1393 1093 1407 1107
rect 1356 927 1363 1073
rect 1376 887 1383 1073
rect 1396 907 1403 1053
rect 1436 987 1443 1113
rect 1456 1087 1463 1216
rect 1376 847 1383 853
rect 1233 833 1247 847
rect 1273 833 1287 847
rect 1313 833 1327 847
rect 1133 813 1147 827
rect 1096 807 1103 813
rect 1036 627 1043 653
rect 1096 647 1103 793
rect 1136 767 1143 813
rect 1236 747 1243 833
rect 1276 767 1283 833
rect 1293 793 1307 807
rect 1296 787 1303 793
rect 1336 723 1343 833
rect 1353 813 1367 827
rect 1373 833 1387 847
rect 1393 813 1407 827
rect 1356 807 1363 813
rect 1396 767 1403 813
rect 1336 716 1363 723
rect 1033 613 1047 627
rect 1116 627 1123 673
rect 1196 667 1203 693
rect 1193 653 1207 667
rect 1153 613 1167 627
rect 1236 647 1243 713
rect 1233 633 1247 647
rect 1016 583 1023 613
rect 1076 607 1083 613
rect 1016 576 1043 583
rect 996 387 1003 413
rect 1036 387 1043 576
rect 1156 547 1163 613
rect 1076 387 1083 493
rect 1116 387 1123 533
rect 993 373 1007 387
rect 1033 383 1047 387
rect 1033 376 1063 383
rect 1033 373 1047 376
rect 1056 327 1063 376
rect 1073 373 1087 387
rect 1093 353 1107 367
rect 1136 367 1143 413
rect 1176 367 1183 393
rect 1216 367 1223 493
rect 1256 387 1263 613
rect 1276 447 1283 673
rect 1316 667 1323 693
rect 1313 653 1327 667
rect 1336 647 1343 693
rect 1356 687 1363 716
rect 1416 647 1423 753
rect 1436 747 1443 913
rect 1436 647 1443 673
rect 1456 667 1463 893
rect 1476 867 1483 1073
rect 1496 987 1503 1093
rect 1516 1083 1523 1153
rect 1556 1127 1563 1253
rect 1576 1247 1583 1573
rect 1596 1507 1603 1573
rect 1636 1567 1643 1576
rect 1653 1573 1667 1576
rect 1676 1567 1683 1573
rect 1673 1553 1687 1567
rect 1713 1563 1727 1567
rect 1736 1563 1743 1773
rect 1776 1767 1783 1793
rect 1796 1763 1803 1793
rect 1816 1787 1823 1793
rect 1856 1787 1863 1816
rect 1873 1813 1887 1816
rect 1833 1773 1847 1787
rect 1893 1783 1907 1787
rect 1916 1783 1923 1973
rect 1936 1827 1943 2033
rect 1893 1776 1923 1783
rect 1893 1773 1907 1776
rect 1836 1767 1843 1773
rect 1796 1756 1823 1763
rect 1776 1743 1783 1753
rect 1776 1736 1803 1743
rect 1796 1607 1803 1736
rect 1816 1607 1823 1756
rect 1836 1627 1843 1713
rect 1773 1573 1787 1587
rect 1793 1593 1807 1607
rect 1813 1583 1827 1587
rect 1836 1583 1843 1593
rect 1813 1576 1843 1583
rect 1813 1573 1827 1576
rect 1713 1556 1743 1563
rect 1713 1553 1727 1556
rect 1616 1327 1623 1513
rect 1653 1313 1667 1327
rect 1633 1293 1647 1307
rect 1576 1147 1583 1173
rect 1533 1083 1547 1087
rect 1516 1076 1547 1083
rect 1533 1073 1547 1076
rect 1573 1073 1587 1087
rect 1536 1007 1543 1073
rect 1576 1047 1583 1073
rect 1536 883 1543 933
rect 1596 887 1603 1293
rect 1616 1147 1623 1193
rect 1636 1187 1643 1293
rect 1656 1287 1663 1313
rect 1676 1147 1683 1353
rect 1696 1347 1703 1473
rect 1736 1347 1743 1393
rect 1756 1347 1763 1553
rect 1776 1547 1783 1573
rect 1796 1487 1803 1553
rect 1836 1407 1843 1553
rect 1856 1547 1863 1653
rect 1936 1627 1943 1813
rect 1976 1744 1984 1856
rect 1956 1627 1963 1633
rect 1953 1613 1967 1627
rect 1893 1573 1907 1587
rect 1933 1573 1947 1587
rect 1973 1573 1987 1587
rect 1896 1567 1903 1573
rect 1693 1333 1707 1347
rect 1713 1313 1727 1327
rect 1733 1333 1747 1347
rect 1696 1267 1703 1293
rect 1716 1287 1723 1313
rect 1833 1293 1847 1307
rect 1696 1147 1703 1153
rect 1636 1107 1643 1133
rect 1676 1107 1683 1113
rect 1633 1093 1647 1107
rect 1673 1093 1687 1107
rect 1696 1087 1703 1133
rect 1693 1073 1707 1087
rect 1616 1067 1623 1073
rect 1616 947 1623 1033
rect 1516 876 1543 883
rect 1516 867 1523 876
rect 1567 876 1573 883
rect 1493 833 1507 847
rect 1513 853 1527 867
rect 1496 787 1503 833
rect 1596 827 1603 853
rect 1476 647 1483 733
rect 1333 633 1347 647
rect 1353 613 1367 627
rect 1433 633 1447 647
rect 1393 623 1407 627
rect 1393 616 1423 623
rect 1393 613 1407 616
rect 1356 527 1363 613
rect 1356 427 1363 433
rect 1376 427 1383 593
rect 1416 587 1423 616
rect 1453 613 1467 627
rect 1473 633 1487 647
rect 1496 627 1503 693
rect 1493 613 1507 627
rect 1456 607 1463 613
rect 1516 547 1523 653
rect 1496 523 1503 533
rect 1536 527 1543 673
rect 1556 647 1563 813
rect 1616 767 1623 913
rect 1636 907 1643 1013
rect 1656 1007 1663 1073
rect 1756 1047 1763 1113
rect 1656 907 1663 933
rect 1633 833 1647 847
rect 1636 827 1643 833
rect 1653 813 1667 827
rect 1693 813 1707 827
rect 1656 707 1663 813
rect 1696 727 1703 813
rect 1716 807 1723 813
rect 1716 703 1723 773
rect 1736 767 1743 873
rect 1756 867 1763 973
rect 1776 947 1783 1193
rect 1796 1147 1803 1273
rect 1836 1267 1843 1293
rect 1856 1227 1863 1393
rect 1916 1367 1923 1573
rect 1936 1387 1943 1573
rect 1893 1333 1907 1347
rect 1873 1313 1887 1327
rect 1876 1307 1883 1313
rect 1856 1107 1863 1133
rect 1876 1127 1883 1293
rect 1896 1287 1903 1333
rect 1916 1123 1923 1313
rect 1936 1267 1943 1293
rect 1956 1267 1963 1573
rect 1976 1567 1983 1573
rect 1996 1567 2003 2013
rect 2016 2007 2023 2053
rect 2076 1947 2083 2056
rect 2113 2053 2127 2067
rect 2153 2053 2167 2067
rect 2173 2073 2187 2087
rect 2196 2063 2203 2196
rect 2216 2127 2223 2273
rect 2235 2224 2243 2304
rect 2256 2287 2263 2353
rect 2276 2247 2283 2313
rect 2296 2267 2303 2633
rect 2336 2287 2343 2513
rect 2356 2307 2363 2773
rect 2416 2767 2423 2976
rect 2436 2787 2443 3036
rect 2456 2987 2463 3013
rect 2476 2807 2483 3013
rect 2496 2827 2503 3573
rect 2536 3547 2543 3693
rect 2555 3664 2563 3744
rect 2616 3707 2623 3973
rect 2676 3967 2683 4233
rect 2713 4173 2727 4187
rect 2753 4173 2767 4187
rect 2716 4087 2723 4173
rect 2756 4127 2763 4173
rect 2796 4144 2804 4256
rect 2816 4087 2823 4476
rect 2833 4473 2847 4476
rect 2895 4436 2903 4516
rect 3147 4516 3163 4523
rect 2913 4483 2927 4487
rect 2936 4483 2943 4493
rect 2913 4476 2943 4483
rect 2913 4473 2927 4476
rect 3016 4427 3023 4513
rect 3056 4487 3063 4513
rect 3096 4487 3103 4513
rect 3156 4507 3163 4516
rect 3176 4507 3183 4513
rect 3153 4493 3167 4507
rect 3053 4473 3067 4487
rect 3093 4473 3107 4487
rect 3116 4467 3123 4493
rect 3136 4487 3143 4493
rect 3133 4473 3147 4487
rect 3176 4487 3183 4493
rect 3236 4487 3243 4513
rect 3336 4507 3343 4533
rect 3333 4493 3347 4507
rect 3173 4473 3187 4487
rect 3233 4473 3247 4487
rect 3213 4463 3227 4467
rect 3196 4456 3227 4463
rect 2895 4398 2903 4422
rect 2916 4147 2923 4213
rect 2993 4173 3007 4187
rect 3033 4173 3047 4187
rect 2996 4147 3003 4173
rect 2696 3924 2704 4036
rect 2736 4007 2743 4033
rect 2733 3993 2747 4007
rect 2835 3956 2843 4036
rect 2893 4023 2907 4027
rect 2853 4003 2867 4007
rect 2876 4016 2907 4023
rect 2876 4003 2883 4016
rect 2853 3996 2883 4003
rect 2893 4013 2907 4016
rect 2956 4007 2963 4133
rect 3036 4127 3043 4173
rect 3076 4167 3083 4433
rect 3116 4267 3123 4433
rect 3196 4427 3203 4456
rect 3213 4453 3227 4456
rect 3313 4483 3327 4487
rect 3296 4476 3327 4483
rect 3296 4467 3303 4476
rect 3313 4473 3327 4476
rect 3376 4463 3383 4473
rect 3376 4456 3393 4463
rect 3196 4227 3203 4273
rect 3133 4223 3147 4227
rect 3133 4216 3163 4223
rect 3133 4213 3147 4216
rect 2996 4007 3003 4033
rect 3056 4007 3063 4013
rect 2953 4003 2967 4007
rect 2853 3993 2867 3996
rect 2573 3703 2587 3707
rect 2573 3696 2603 3703
rect 2573 3693 2587 3696
rect 2596 3667 2603 3696
rect 2653 3693 2667 3707
rect 2733 3723 2747 3727
rect 2716 3716 2747 3723
rect 2716 3707 2723 3716
rect 2733 3713 2747 3716
rect 2693 3703 2707 3707
rect 2693 3696 2713 3703
rect 2693 3693 2707 3696
rect 2656 3687 2663 3693
rect 2536 3527 2543 3533
rect 2576 3527 2583 3553
rect 2533 3523 2547 3527
rect 2533 3516 2563 3523
rect 2533 3513 2547 3516
rect 2516 3127 2523 3353
rect 2533 3223 2547 3227
rect 2556 3223 2563 3516
rect 2573 3513 2587 3527
rect 2616 3444 2624 3556
rect 2676 3527 2683 3673
rect 2756 3667 2763 3673
rect 2776 3627 2783 3953
rect 2835 3918 2843 3942
rect 2793 3693 2807 3707
rect 2833 3703 2847 3707
rect 2856 3703 2863 3993
rect 2936 3996 2967 4003
rect 2936 3967 2943 3996
rect 2953 3993 2967 3996
rect 2993 3993 3007 4007
rect 3053 3993 3067 4007
rect 3096 4007 3103 4153
rect 3156 4127 3163 4216
rect 3193 4213 3207 4227
rect 3213 4193 3227 4207
rect 3216 4187 3223 4193
rect 3256 4167 3263 4253
rect 3276 4227 3283 4233
rect 3273 4213 3287 4227
rect 3333 4173 3347 4187
rect 3336 4167 3343 4173
rect 3373 4173 3387 4187
rect 3376 4167 3383 4173
rect 3353 4153 3367 4167
rect 3356 4067 3363 4153
rect 2796 3687 2803 3693
rect 2833 3696 2863 3703
rect 2833 3693 2847 3696
rect 2813 3673 2827 3687
rect 2816 3647 2823 3673
rect 2716 3527 2723 3553
rect 2713 3513 2727 3527
rect 2773 3523 2787 3527
rect 2756 3516 2787 3523
rect 2533 3216 2563 3223
rect 2533 3213 2547 3216
rect 2556 3207 2563 3216
rect 2573 3213 2587 3227
rect 2516 3047 2523 3113
rect 2553 3043 2567 3047
rect 2576 3043 2583 3213
rect 2616 3184 2624 3296
rect 2673 3213 2687 3227
rect 2676 3167 2683 3213
rect 2616 3047 2623 3053
rect 2553 3036 2583 3043
rect 2553 3033 2567 3036
rect 2613 3033 2627 3047
rect 2573 3023 2587 3027
rect 2573 3016 2603 3023
rect 2573 3013 2587 3016
rect 2476 2767 2483 2773
rect 2376 2607 2383 2753
rect 2393 2733 2407 2747
rect 2396 2647 2403 2733
rect 2473 2753 2487 2767
rect 2413 2713 2427 2727
rect 2453 2713 2467 2727
rect 2416 2583 2423 2713
rect 2456 2707 2463 2713
rect 2416 2576 2443 2583
rect 2436 2567 2443 2576
rect 2496 2583 2503 2793
rect 2536 2723 2543 2993
rect 2596 2987 2603 3016
rect 2636 2807 2643 3133
rect 2696 3047 2703 3493
rect 2756 3427 2763 3516
rect 2773 3513 2787 3516
rect 2836 3483 2843 3513
rect 2853 3483 2867 3487
rect 2836 3476 2867 3483
rect 2853 3473 2867 3476
rect 2713 3213 2727 3227
rect 2716 3187 2723 3213
rect 2716 3107 2723 3173
rect 2756 3067 2763 3413
rect 2797 3278 2805 3302
rect 2797 3184 2805 3264
rect 2853 3213 2867 3227
rect 2893 3213 2907 3227
rect 2676 3003 2683 3033
rect 2693 3003 2707 3007
rect 2676 2996 2707 3003
rect 2693 2993 2707 2996
rect 2596 2743 2603 2773
rect 2613 2743 2627 2747
rect 2596 2736 2627 2743
rect 2673 2763 2687 2767
rect 2696 2763 2703 2993
rect 2776 2867 2783 3153
rect 2673 2756 2703 2763
rect 2673 2753 2687 2756
rect 2613 2733 2627 2736
rect 2653 2733 2667 2747
rect 2713 2733 2727 2747
rect 2516 2716 2543 2723
rect 2516 2667 2523 2716
rect 2496 2576 2523 2583
rect 2433 2563 2447 2567
rect 2453 2563 2467 2567
rect 2433 2556 2467 2563
rect 2433 2553 2447 2556
rect 2453 2553 2467 2556
rect 2516 2347 2523 2576
rect 2536 2567 2543 2693
rect 2533 2553 2547 2567
rect 2556 2507 2563 2733
rect 2656 2727 2663 2733
rect 2716 2727 2723 2733
rect 2796 2707 2803 3053
rect 2816 2964 2824 3076
rect 2836 3007 2843 3213
rect 2856 3207 2863 3213
rect 2856 3107 2863 3193
rect 2896 3167 2903 3213
rect 2856 3047 2863 3073
rect 2853 3033 2867 3047
rect 2816 2787 2823 2793
rect 2813 2773 2827 2787
rect 2876 2727 2883 3093
rect 2896 3047 2903 3093
rect 2893 3033 2907 3047
rect 2916 2787 2923 3613
rect 2936 3527 2943 3953
rect 2976 3727 2983 3973
rect 3173 3953 3187 3967
rect 3176 3947 3183 3953
rect 3156 3727 3163 3753
rect 3216 3743 3223 4013
rect 3236 4007 3243 4033
rect 3233 3993 3247 4007
rect 3316 4007 3323 4013
rect 3293 3973 3307 3987
rect 3313 3993 3327 4007
rect 3216 3736 3243 3743
rect 3033 3723 3047 3727
rect 3093 3723 3107 3727
rect 2953 3693 2967 3707
rect 2956 3687 2963 3693
rect 2993 3693 3007 3707
rect 3033 3716 3063 3723
rect 3033 3713 3047 3716
rect 2973 3673 2987 3687
rect 2956 3667 2963 3673
rect 2976 3623 2983 3673
rect 2996 3647 3003 3693
rect 3013 3673 3027 3687
rect 3016 3623 3023 3673
rect 2976 3616 3023 3623
rect 3056 3607 3063 3716
rect 3076 3716 3107 3723
rect 3076 3687 3083 3716
rect 3093 3713 3107 3716
rect 3133 3693 3147 3707
rect 3193 3713 3207 3727
rect 3173 3693 3187 3707
rect 3113 3673 3127 3687
rect 3116 3667 3123 3673
rect 3136 3647 3143 3693
rect 3176 3587 3183 3693
rect 3196 3687 3203 3713
rect 3216 3567 3223 3713
rect 2953 3513 2967 3527
rect 2956 3487 2963 3513
rect 2977 3476 2985 3556
rect 3036 3527 3043 3533
rect 3033 3513 3047 3527
rect 2936 3184 2944 3296
rect 2956 3247 2963 3473
rect 2977 3438 2985 3462
rect 2976 3127 2983 3213
rect 2955 2996 2963 3076
rect 2973 3033 2987 3047
rect 2976 2987 2983 3033
rect 2996 3007 3003 3453
rect 3116 3444 3124 3556
rect 3236 3547 3243 3736
rect 3276 3727 3283 3733
rect 3296 3727 3303 3973
rect 3336 3727 3343 4013
rect 3356 4007 3363 4053
rect 3376 3727 3383 3953
rect 3396 3747 3403 4233
rect 3436 4167 3443 4533
rect 3477 4436 3485 4516
rect 3477 4398 3485 4422
rect 3456 4144 3464 4256
rect 3496 4247 3503 4513
rect 3533 4483 3547 4487
rect 3516 4476 3547 4483
rect 3516 4183 3523 4476
rect 3533 4473 3547 4476
rect 3616 4404 3624 4516
rect 3595 4238 3603 4262
rect 3533 4183 3547 4187
rect 3516 4176 3547 4183
rect 3533 4173 3547 4176
rect 3536 4087 3543 4173
rect 3595 4144 3603 4224
rect 3616 4187 3623 4213
rect 3533 4023 3547 4027
rect 3556 4023 3563 4093
rect 3533 4016 3563 4023
rect 3533 4013 3547 4016
rect 3476 4007 3483 4013
rect 3373 3713 3387 3727
rect 3293 3673 3307 3687
rect 3393 3693 3407 3707
rect 3353 3673 3367 3687
rect 3296 3627 3303 3673
rect 3356 3667 3363 3673
rect 3096 3247 3103 3273
rect 3136 3267 3143 3513
rect 3156 3327 3163 3533
rect 3216 3527 3223 3533
rect 3213 3513 3227 3527
rect 3176 3487 3183 3513
rect 3236 3467 3243 3493
rect 3276 3307 3283 3553
rect 3356 3547 3363 3553
rect 3353 3533 3367 3547
rect 3336 3527 3343 3533
rect 3293 3493 3307 3507
rect 3333 3513 3347 3527
rect 3376 3527 3383 3673
rect 3396 3647 3403 3693
rect 3416 3627 3423 3993
rect 3473 3993 3487 4007
rect 3573 3993 3587 4007
rect 3576 3947 3583 3993
rect 3597 3956 3605 4036
rect 3597 3918 3605 3942
rect 3636 3927 3643 4493
rect 3673 4483 3687 4487
rect 3656 4476 3687 4483
rect 3656 4447 3663 4476
rect 3673 4473 3687 4476
rect 3873 4453 3887 4467
rect 3813 4433 3827 4447
rect 3656 4167 3663 4233
rect 3716 4227 3723 4233
rect 3693 4193 3707 4207
rect 3713 4213 3727 4227
rect 3696 4107 3703 4193
rect 3733 4173 3747 4187
rect 3736 4167 3743 4173
rect 3753 4153 3767 4167
rect 3656 4007 3663 4073
rect 3653 3993 3667 4007
rect 3676 3967 3683 4033
rect 3736 3924 3744 4036
rect 3756 4027 3763 4153
rect 3776 3907 3783 4153
rect 3453 3723 3467 3727
rect 3453 3716 3483 3723
rect 3453 3713 3467 3716
rect 3396 3547 3403 3553
rect 3436 3547 3443 3613
rect 3373 3523 3387 3527
rect 3373 3516 3403 3523
rect 3373 3513 3387 3516
rect 3396 3507 3403 3516
rect 3296 3487 3303 3493
rect 3296 3283 3303 3393
rect 3276 3276 3303 3283
rect 3216 3247 3223 3273
rect 3113 3233 3127 3247
rect 3073 3213 3087 3227
rect 3036 3047 3043 3193
rect 3076 3187 3083 3213
rect 3096 3207 3103 3233
rect 3116 3227 3123 3233
rect 3173 3213 3187 3227
rect 3193 3213 3207 3227
rect 3213 3233 3227 3247
rect 3253 3233 3267 3247
rect 3176 3207 3183 3213
rect 3076 3047 3083 3173
rect 2955 2958 2963 2982
rect 2636 2567 2643 2673
rect 2593 2563 2607 2567
rect 2593 2556 2623 2563
rect 2593 2553 2607 2556
rect 2333 2273 2347 2287
rect 2213 2063 2227 2067
rect 2196 2056 2227 2063
rect 2156 1947 2163 2053
rect 2013 1773 2027 1787
rect 2053 1783 2067 1787
rect 2076 1783 2083 1813
rect 2053 1776 2083 1783
rect 2053 1773 2067 1776
rect 2016 1627 2023 1773
rect 2036 1607 2043 1633
rect 2096 1607 2103 1933
rect 2196 1867 2203 2056
rect 2213 2053 2227 2056
rect 2236 1987 2243 2153
rect 2115 1838 2123 1862
rect 2115 1744 2123 1824
rect 2156 1647 2163 1833
rect 2196 1827 2203 1853
rect 2256 1807 2263 2213
rect 2276 1847 2283 2093
rect 2176 1627 2183 1793
rect 2196 1623 2203 1773
rect 2233 1773 2247 1787
rect 2236 1763 2243 1773
rect 2253 1763 2267 1767
rect 2236 1756 2283 1763
rect 2253 1753 2267 1756
rect 2213 1623 2227 1627
rect 2196 1616 2227 1623
rect 2213 1613 2227 1616
rect 2156 1607 2163 1613
rect 2153 1593 2167 1607
rect 2016 1587 2023 1593
rect 2013 1573 2027 1587
rect 2096 1567 2103 1593
rect 2136 1587 2143 1593
rect 2133 1573 2147 1587
rect 2173 1573 2187 1587
rect 2276 1603 2283 1756
rect 2296 1727 2303 2133
rect 2353 2053 2367 2067
rect 2336 1827 2343 2053
rect 2356 1847 2363 2053
rect 2376 1987 2383 2233
rect 2396 2107 2403 2293
rect 2493 2273 2507 2287
rect 2453 2243 2467 2247
rect 2496 2243 2503 2273
rect 2536 2247 2543 2273
rect 2576 2267 2583 2493
rect 2616 2327 2623 2556
rect 2633 2553 2647 2567
rect 2653 2533 2667 2547
rect 2696 2547 2703 2593
rect 2656 2507 2663 2533
rect 2716 2507 2723 2693
rect 2813 2583 2827 2587
rect 2796 2576 2827 2583
rect 2796 2567 2803 2576
rect 2813 2573 2827 2576
rect 2836 2567 2843 2573
rect 2833 2553 2847 2567
rect 2736 2523 2743 2553
rect 2753 2523 2767 2527
rect 2736 2516 2767 2523
rect 2856 2527 2863 2573
rect 2873 2533 2887 2547
rect 2753 2513 2767 2516
rect 2876 2507 2883 2533
rect 2636 2307 2643 2353
rect 2633 2293 2647 2307
rect 2593 2263 2607 2267
rect 2616 2263 2623 2293
rect 2593 2256 2623 2263
rect 2593 2253 2607 2256
rect 2653 2253 2667 2267
rect 2453 2236 2503 2243
rect 2453 2233 2467 2236
rect 2393 2033 2407 2047
rect 2433 2043 2447 2047
rect 2456 2043 2463 2193
rect 2496 2087 2503 2236
rect 2493 2073 2507 2087
rect 2433 2036 2463 2043
rect 2433 2033 2447 2036
rect 2513 2033 2527 2047
rect 2396 1947 2403 2033
rect 2516 1967 2523 2033
rect 2313 1773 2327 1787
rect 2353 1773 2367 1787
rect 2316 1763 2323 1773
rect 2316 1756 2343 1763
rect 2293 1603 2307 1607
rect 2276 1596 2307 1603
rect 2293 1593 2307 1596
rect 2073 1553 2087 1567
rect 2076 1543 2083 1553
rect 2116 1547 2123 1573
rect 2176 1567 2183 1573
rect 2317 1556 2325 1636
rect 2336 1567 2343 1756
rect 2356 1747 2363 1773
rect 2076 1536 2093 1543
rect 1996 1347 2003 1533
rect 2317 1518 2325 1542
rect 1973 1293 1987 1307
rect 2013 1293 2027 1307
rect 1976 1287 1983 1293
rect 1916 1116 1943 1123
rect 1793 1073 1807 1087
rect 1833 1073 1847 1087
rect 1853 1093 1867 1107
rect 1796 1067 1803 1073
rect 1836 1067 1843 1073
rect 1936 1067 1943 1116
rect 1976 1107 1983 1273
rect 2016 1247 2023 1293
rect 1953 1073 1967 1087
rect 1973 1093 1987 1107
rect 1993 1073 2007 1087
rect 1756 747 1763 813
rect 1796 807 1803 973
rect 1816 967 1823 1033
rect 1816 827 1823 953
rect 1836 927 1843 1053
rect 1956 1047 1963 1073
rect 1996 1063 2003 1073
rect 1976 1056 2003 1063
rect 1836 847 1843 873
rect 1896 867 1903 1013
rect 1936 887 1943 893
rect 1936 867 1943 873
rect 1976 867 1983 1056
rect 2016 1027 2023 1213
rect 2056 1147 2063 1373
rect 2096 1327 2103 1373
rect 2356 1347 2363 1633
rect 2373 1603 2387 1607
rect 2396 1603 2403 1853
rect 2413 1773 2427 1787
rect 2416 1767 2423 1773
rect 2453 1773 2467 1787
rect 2433 1753 2447 1767
rect 2416 1607 2423 1733
rect 2436 1647 2443 1753
rect 2456 1747 2463 1773
rect 2476 1743 2483 1833
rect 2536 1823 2543 2153
rect 2596 2087 2603 2153
rect 2593 2073 2607 2087
rect 2616 2007 2623 2233
rect 2656 2227 2663 2253
rect 2676 2167 2683 2333
rect 2737 2318 2745 2342
rect 2713 2263 2727 2267
rect 2696 2256 2727 2263
rect 2696 2207 2703 2256
rect 2713 2253 2727 2256
rect 2737 2224 2745 2304
rect 2633 2063 2647 2067
rect 2656 2063 2663 2133
rect 2633 2056 2663 2063
rect 2633 2053 2647 2056
rect 2676 2047 2683 2073
rect 2693 2033 2707 2047
rect 2696 2007 2703 2033
rect 2536 1816 2563 1823
rect 2496 1767 2503 1773
rect 2513 1753 2527 1767
rect 2516 1747 2523 1753
rect 2476 1736 2503 1743
rect 2373 1596 2403 1603
rect 2373 1593 2387 1596
rect 2413 1593 2427 1607
rect 2153 1333 2167 1347
rect 2156 1327 2163 1333
rect 2093 1313 2107 1327
rect 2133 1313 2147 1327
rect 2233 1343 2247 1347
rect 2216 1336 2247 1343
rect 2136 1287 2143 1313
rect 2096 1127 2103 1253
rect 2136 1127 2143 1233
rect 2053 1123 2067 1127
rect 2036 1116 2067 1123
rect 2036 1067 2043 1116
rect 2053 1113 2067 1116
rect 2073 1093 2087 1107
rect 2093 1113 2107 1127
rect 2156 1107 2163 1293
rect 2216 1247 2223 1336
rect 2233 1333 2247 1336
rect 2253 1313 2267 1327
rect 2376 1327 2383 1533
rect 2436 1363 2443 1613
rect 2456 1524 2464 1636
rect 2416 1356 2443 1363
rect 2256 1307 2263 1313
rect 2373 1313 2387 1327
rect 2313 1283 2327 1287
rect 2296 1276 2327 1283
rect 2216 1127 2223 1133
rect 2076 1087 2083 1093
rect 2216 1087 2223 1113
rect 2296 1107 2303 1276
rect 2313 1273 2327 1276
rect 2233 1103 2247 1107
rect 2233 1096 2263 1103
rect 2233 1093 2247 1096
rect 2213 1073 2227 1087
rect 2256 1067 2263 1096
rect 2293 1093 2307 1107
rect 2333 1093 2347 1107
rect 2313 1083 2327 1087
rect 2336 1083 2343 1093
rect 2313 1076 2343 1083
rect 2313 1073 2327 1076
rect 2316 1067 2323 1073
rect 1893 853 1907 867
rect 1833 833 1847 847
rect 1853 793 1867 807
rect 1856 787 1863 793
rect 1696 696 1723 703
rect 1596 667 1603 673
rect 1553 633 1567 647
rect 1573 613 1587 627
rect 1613 623 1627 627
rect 1696 647 1703 696
rect 1633 623 1647 627
rect 1613 616 1647 623
rect 1613 613 1627 616
rect 1633 613 1647 616
rect 1673 613 1687 627
rect 1693 633 1707 647
rect 1576 607 1583 613
rect 1496 516 1523 523
rect 1276 367 1283 373
rect 956 167 963 193
rect 996 187 1003 313
rect 1016 187 1023 213
rect 1036 207 1043 293
rect 1096 227 1103 353
rect 1173 353 1187 367
rect 1193 333 1207 347
rect 1213 353 1227 367
rect 1273 353 1287 367
rect 1293 333 1307 347
rect 1116 227 1123 313
rect 1013 173 1027 187
rect 893 133 907 147
rect 953 153 967 167
rect 976 147 983 173
rect 1036 167 1043 193
rect 1076 167 1083 193
rect 1096 167 1103 213
rect 1136 167 1143 293
rect 1176 167 1183 313
rect 1196 287 1203 333
rect 1256 307 1263 333
rect 993 133 1007 147
rect 1033 153 1047 167
rect 1073 153 1087 167
rect 1133 153 1147 167
rect 1096 147 1103 153
rect 1093 133 1107 147
rect 1153 133 1167 147
rect 1173 153 1187 167
rect 996 127 1003 133
rect 1116 123 1123 133
rect 1156 123 1163 133
rect 1116 116 1163 123
rect 976 87 983 113
rect 1216 67 1223 193
rect 1276 147 1283 233
rect 1296 207 1303 333
rect 1336 287 1343 373
rect 1356 367 1363 413
rect 1396 367 1403 453
rect 1456 367 1463 393
rect 1373 333 1387 347
rect 1376 267 1383 333
rect 1433 333 1447 347
rect 1453 353 1467 367
rect 1493 353 1507 367
rect 1393 313 1407 327
rect 1396 267 1403 313
rect 1416 247 1423 313
rect 1436 287 1443 333
rect 1273 133 1287 147
rect 1316 27 1323 173
rect 1336 147 1343 153
rect 1376 147 1383 233
rect 1436 167 1443 173
rect 1456 167 1463 313
rect 1476 267 1483 313
rect 1496 307 1503 353
rect 1516 187 1523 516
rect 1536 367 1543 513
rect 1556 387 1563 513
rect 1576 387 1583 593
rect 1596 527 1603 613
rect 1636 527 1643 613
rect 1676 603 1683 613
rect 1716 607 1723 653
rect 1736 627 1743 673
rect 1776 627 1783 653
rect 1733 623 1747 627
rect 1733 616 1753 623
rect 1733 613 1747 616
rect 1773 613 1787 627
rect 1676 596 1703 603
rect 1553 363 1567 367
rect 1553 356 1583 363
rect 1553 353 1567 356
rect 1533 313 1547 327
rect 1536 287 1543 313
rect 1576 267 1583 356
rect 1596 287 1603 433
rect 1656 407 1663 533
rect 1636 367 1643 393
rect 1676 387 1683 573
rect 1696 527 1703 596
rect 1793 593 1807 607
rect 1716 463 1723 473
rect 1696 456 1723 463
rect 1696 427 1703 456
rect 1716 367 1723 413
rect 1736 367 1743 493
rect 1776 487 1783 573
rect 1796 487 1803 593
rect 1816 547 1823 653
rect 1836 647 1843 753
rect 1876 687 1883 853
rect 1913 833 1927 847
rect 1933 853 1947 867
rect 1976 847 1983 853
rect 1973 833 1987 847
rect 1916 807 1923 833
rect 1833 633 1847 647
rect 1873 643 1887 647
rect 1853 613 1867 627
rect 1873 636 1893 643
rect 1873 633 1887 636
rect 1893 623 1907 627
rect 1893 616 1923 623
rect 1893 613 1907 616
rect 1836 527 1843 593
rect 1856 587 1863 613
rect 1896 567 1903 573
rect 1816 387 1823 393
rect 1773 373 1787 387
rect 1613 333 1627 347
rect 1616 207 1623 333
rect 1653 313 1667 327
rect 1656 267 1663 313
rect 1676 243 1683 313
rect 1696 307 1703 313
rect 1736 283 1743 333
rect 1756 307 1763 333
rect 1736 276 1763 283
rect 1656 236 1683 243
rect 1453 153 1467 167
rect 1436 147 1443 153
rect 1333 133 1347 147
rect 1373 133 1387 147
rect 1536 147 1543 193
rect 1513 133 1527 147
rect 1516 127 1523 133
rect 1393 113 1407 127
rect 1556 127 1563 153
rect 1616 147 1623 193
rect 1553 113 1567 127
rect 1636 127 1643 233
rect 1656 167 1663 236
rect 1696 203 1703 233
rect 1676 196 1703 203
rect 1676 187 1683 196
rect 1653 153 1667 167
rect 1736 147 1743 173
rect 1756 167 1763 276
rect 1776 267 1783 373
rect 1793 353 1807 367
rect 1813 373 1827 387
rect 1796 287 1803 353
rect 1836 347 1843 493
rect 1916 467 1923 616
rect 1856 367 1863 433
rect 1876 367 1883 453
rect 1896 367 1903 413
rect 1916 407 1923 433
rect 1936 403 1943 773
rect 1956 727 1963 793
rect 1996 787 2003 873
rect 2036 867 2043 1053
rect 2033 853 2047 867
rect 2073 853 2087 867
rect 1976 703 1983 733
rect 1956 696 1983 703
rect 1956 647 1963 696
rect 1996 667 2003 753
rect 2016 667 2023 793
rect 1993 653 2007 667
rect 1953 633 1967 647
rect 2036 647 2043 713
rect 2056 707 2063 773
rect 2076 647 2083 853
rect 2093 833 2107 847
rect 2096 803 2103 833
rect 2113 803 2127 807
rect 2096 796 2127 803
rect 2113 793 2127 796
rect 1973 613 1987 627
rect 2013 613 2027 627
rect 2033 633 2047 647
rect 2053 613 2067 627
rect 2073 633 2087 647
rect 2096 627 2103 693
rect 2116 667 2123 793
rect 1976 607 1983 613
rect 1996 487 2003 613
rect 2016 563 2023 613
rect 2016 556 2043 563
rect 2036 547 2043 556
rect 1936 396 1953 403
rect 1956 387 1963 393
rect 2016 387 2023 533
rect 2056 527 2063 613
rect 2116 607 2123 633
rect 2036 387 2043 413
rect 2096 407 2103 553
rect 2116 427 2123 573
rect 2136 527 2143 733
rect 2156 687 2163 933
rect 2233 833 2247 847
rect 2236 807 2243 833
rect 2276 827 2283 1053
rect 2416 887 2423 1356
rect 2476 1347 2483 1673
rect 2496 1507 2503 1736
rect 2536 1607 2543 1773
rect 2556 1687 2563 1816
rect 2573 1773 2587 1787
rect 2613 1783 2627 1787
rect 2656 1783 2663 1973
rect 2613 1776 2663 1783
rect 2676 1823 2683 1953
rect 2736 1847 2743 2033
rect 2693 1823 2707 1827
rect 2676 1816 2707 1823
rect 2613 1773 2627 1776
rect 2576 1767 2583 1773
rect 2556 1607 2563 1653
rect 2676 1647 2683 1816
rect 2693 1813 2707 1816
rect 2713 1793 2727 1807
rect 2716 1783 2723 1793
rect 2707 1776 2723 1783
rect 2756 1647 2763 1993
rect 2816 1947 2823 2493
rect 2833 2263 2847 2267
rect 2856 2263 2863 2273
rect 2833 2256 2863 2263
rect 2833 2253 2847 2256
rect 2876 2224 2884 2336
rect 2896 2187 2903 2573
rect 2916 2567 2923 2773
rect 2936 2704 2944 2816
rect 2956 2563 2963 2833
rect 2996 2647 3003 2853
rect 3013 2733 3027 2747
rect 3016 2727 3023 2733
rect 3036 2687 3043 2993
rect 2996 2567 3003 2633
rect 3036 2567 3043 2573
rect 2956 2556 2983 2563
rect 2953 2513 2967 2527
rect 2956 2507 2963 2513
rect 2976 2427 2983 2556
rect 2993 2553 3007 2567
rect 3033 2553 3047 2567
rect 2916 2167 2923 2413
rect 3056 2323 3063 2973
rect 3096 2947 3103 3053
rect 3116 3047 3123 3073
rect 3156 3067 3163 3073
rect 3153 3053 3167 3067
rect 3113 3033 3127 3047
rect 3196 3047 3203 3213
rect 3256 3127 3263 3233
rect 3276 3207 3283 3276
rect 3416 3247 3423 3473
rect 3456 3283 3463 3653
rect 3476 3567 3483 3716
rect 3493 3703 3507 3707
rect 3516 3703 3523 3753
rect 3493 3696 3523 3703
rect 3493 3693 3507 3696
rect 3576 3703 3583 3733
rect 3616 3727 3623 3753
rect 3593 3703 3607 3707
rect 3576 3696 3607 3703
rect 3613 3713 3627 3727
rect 3653 3723 3667 3727
rect 3676 3723 3683 3833
rect 3653 3716 3683 3723
rect 3653 3713 3667 3716
rect 3633 3703 3647 3707
rect 3693 3703 3707 3707
rect 3593 3693 3607 3696
rect 3633 3696 3707 3703
rect 3753 3713 3767 3727
rect 3633 3693 3647 3696
rect 3693 3693 3707 3696
rect 3596 3607 3603 3693
rect 3476 3347 3483 3533
rect 3496 3527 3503 3593
rect 3493 3513 3507 3527
rect 3536 3527 3543 3553
rect 3576 3547 3583 3553
rect 3573 3533 3587 3547
rect 3533 3513 3547 3527
rect 3593 3493 3607 3507
rect 3436 3276 3463 3283
rect 3436 3267 3443 3276
rect 3313 3233 3327 3247
rect 3133 3013 3147 3027
rect 3233 3043 3247 3047
rect 3233 3036 3263 3043
rect 3233 3033 3247 3036
rect 3136 3007 3143 3013
rect 3096 2887 3103 2933
rect 3075 2798 3083 2822
rect 3075 2704 3083 2784
rect 3096 2747 3103 2793
rect 3093 2733 3107 2747
rect 3116 2567 3123 2693
rect 3156 2667 3163 3013
rect 3256 2987 3263 3036
rect 3176 2704 3184 2816
rect 3213 2733 3227 2747
rect 3253 2733 3267 2747
rect 3216 2707 3223 2733
rect 3256 2727 3263 2733
rect 3276 2703 3283 3193
rect 3296 3007 3303 3233
rect 3316 3227 3323 3233
rect 3333 3213 3347 3227
rect 3393 3213 3407 3227
rect 3413 3233 3427 3247
rect 3453 3233 3467 3247
rect 3456 3227 3463 3233
rect 3433 3213 3447 3227
rect 3336 3167 3343 3213
rect 3376 3087 3383 3213
rect 3396 3207 3403 3213
rect 3256 2696 3283 2703
rect 3113 2553 3127 2567
rect 3036 2316 3063 2323
rect 2996 2287 3003 2293
rect 2953 2273 2967 2287
rect 2936 2247 2943 2253
rect 2876 2004 2884 2116
rect 2936 2083 2943 2233
rect 2956 2207 2963 2273
rect 2993 2273 3007 2287
rect 3013 2253 3027 2267
rect 3016 2187 3023 2253
rect 2953 2083 2967 2087
rect 2936 2076 2967 2083
rect 2776 1687 2783 1773
rect 2813 1773 2827 1787
rect 2833 1773 2847 1787
rect 2916 1787 2923 2033
rect 2936 1867 2943 2076
rect 2953 2073 2967 2076
rect 2816 1767 2823 1773
rect 2836 1767 2843 1773
rect 2933 1753 2947 1767
rect 2596 1607 2603 1613
rect 2553 1593 2567 1607
rect 2593 1593 2607 1607
rect 2616 1567 2623 1633
rect 2716 1607 2723 1633
rect 2796 1623 2803 1753
rect 2836 1627 2843 1673
rect 2936 1647 2943 1753
rect 2813 1623 2827 1627
rect 2796 1616 2827 1623
rect 2713 1593 2727 1607
rect 2813 1613 2827 1616
rect 2767 1596 2783 1603
rect 2776 1567 2783 1596
rect 2453 1313 2467 1327
rect 2456 1287 2463 1313
rect 2556 1303 2563 1553
rect 2796 1547 2803 1573
rect 2596 1307 2603 1333
rect 2656 1327 2663 1353
rect 2573 1303 2587 1307
rect 2556 1296 2587 1303
rect 2573 1293 2587 1296
rect 2613 1293 2627 1307
rect 2653 1313 2667 1327
rect 2693 1323 2707 1327
rect 2716 1323 2723 1333
rect 2816 1327 2823 1333
rect 2693 1316 2723 1323
rect 2693 1313 2707 1316
rect 2793 1293 2807 1307
rect 2616 1147 2623 1293
rect 2796 1247 2803 1293
rect 2473 1143 2487 1147
rect 2473 1136 2503 1143
rect 2473 1133 2487 1136
rect 2496 967 2503 1136
rect 2636 1127 2643 1173
rect 2676 1127 2683 1153
rect 2696 1147 2703 1193
rect 2696 1127 2703 1133
rect 2633 1113 2647 1127
rect 2673 1113 2687 1127
rect 2693 1113 2707 1127
rect 2656 1087 2663 1093
rect 2356 847 2363 853
rect 2453 853 2467 867
rect 2293 813 2307 827
rect 2353 833 2367 847
rect 2296 807 2303 813
rect 2333 793 2347 807
rect 2373 793 2387 807
rect 2176 627 2183 793
rect 2196 607 2203 753
rect 2236 647 2243 673
rect 2256 647 2263 773
rect 2276 647 2283 733
rect 2336 687 2343 793
rect 2376 707 2383 793
rect 2316 647 2323 653
rect 2336 647 2343 653
rect 2376 647 2383 673
rect 2273 633 2287 647
rect 2216 627 2223 633
rect 2213 623 2227 627
rect 2253 623 2267 627
rect 2213 616 2267 623
rect 2213 613 2227 616
rect 2176 547 2183 573
rect 2136 403 2143 473
rect 2176 407 2183 473
rect 2116 396 2143 403
rect 2116 387 2123 396
rect 1953 373 1967 387
rect 1853 353 1867 367
rect 1893 353 1907 367
rect 1776 147 1783 193
rect 1713 133 1727 147
rect 1396 107 1403 113
rect 1476 -24 1483 73
rect 1516 67 1523 113
rect 1696 107 1703 133
rect 1716 127 1723 133
rect 1773 133 1787 147
rect 1816 127 1823 333
rect 1873 313 1887 327
rect 1856 147 1863 313
rect 1876 267 1883 313
rect 1793 113 1807 127
rect 1833 113 1847 127
rect 1853 133 1867 147
rect 1873 113 1887 127
rect 1796 107 1803 113
rect 1836 87 1843 113
rect 1756 -24 1763 53
rect 1876 47 1883 113
rect 1896 -24 1903 113
rect 1916 87 1923 113
rect 1936 47 1943 373
rect 1973 353 1987 367
rect 2033 373 2047 387
rect 2113 373 2127 387
rect 2153 383 2167 387
rect 1956 187 1963 293
rect 1976 267 1983 353
rect 2016 327 2023 353
rect 2096 343 2103 373
rect 2153 376 2183 383
rect 2153 373 2167 376
rect 2096 336 2123 343
rect 2036 307 2043 313
rect 1956 167 1963 173
rect 1953 153 1967 167
rect 1936 -24 1943 33
rect 1976 27 1983 153
rect 1996 107 2003 293
rect 2016 167 2023 213
rect 2056 187 2063 333
rect 2076 187 2083 233
rect 2096 207 2103 313
rect 2033 123 2047 127
rect 2056 123 2063 173
rect 2076 167 2083 173
rect 2096 167 2103 193
rect 2073 153 2087 167
rect 2093 153 2107 167
rect 2033 116 2063 123
rect 2033 113 2047 116
rect 2056 87 2063 116
rect 2116 67 2123 336
rect 2136 307 2143 353
rect 2176 227 2183 376
rect 2196 367 2203 453
rect 2216 387 2223 553
rect 2236 367 2243 616
rect 2253 613 2267 616
rect 2313 633 2327 647
rect 2333 633 2347 647
rect 2373 633 2387 647
rect 2396 627 2403 633
rect 2393 613 2407 627
rect 2276 447 2283 593
rect 2296 487 2303 593
rect 2416 507 2423 653
rect 2436 627 2443 753
rect 2456 707 2463 853
rect 2473 833 2487 847
rect 2476 687 2483 833
rect 2516 667 2523 973
rect 2556 867 2563 953
rect 2796 867 2803 1113
rect 2816 1044 2824 1156
rect 2856 1127 2863 1173
rect 2876 1167 2883 1573
rect 2896 1567 2903 1593
rect 2896 1264 2904 1376
rect 2896 1127 2903 1153
rect 2853 1113 2867 1127
rect 2893 1113 2907 1127
rect 2916 1067 2923 1533
rect 2976 1367 2983 2173
rect 3036 2127 3043 2316
rect 3096 2287 3103 2353
rect 3156 2307 3163 2653
rect 3156 2287 3163 2293
rect 3053 2273 3067 2287
rect 3056 2267 3063 2273
rect 3093 2273 3107 2287
rect 3113 2253 3127 2267
rect 3133 2253 3147 2267
rect 3153 2273 3167 2287
rect 3193 2273 3207 2287
rect 3196 2267 3203 2273
rect 3116 2207 3123 2253
rect 2996 1627 3003 2113
rect 3015 2036 3023 2116
rect 3116 2103 3123 2193
rect 3136 2187 3143 2253
rect 3216 2227 3223 2673
rect 3236 2567 3243 2593
rect 3233 2553 3247 2567
rect 3256 2467 3263 2696
rect 3296 2627 3303 2993
rect 3316 2964 3324 3076
rect 3396 3047 3403 3093
rect 3436 3047 3443 3213
rect 3476 3207 3483 3313
rect 3496 3267 3503 3473
rect 3536 3267 3543 3333
rect 3493 3253 3507 3267
rect 3513 3233 3527 3247
rect 3393 3033 3407 3047
rect 3455 2996 3463 3076
rect 3473 3043 3487 3047
rect 3496 3043 3503 3073
rect 3473 3036 3503 3043
rect 3473 3033 3487 3036
rect 3315 2798 3323 2822
rect 3315 2704 3323 2784
rect 3333 2743 3347 2747
rect 3333 2736 3363 2743
rect 3333 2733 3347 2736
rect 3356 2587 3363 2736
rect 3336 2567 3343 2573
rect 3376 2567 3383 2953
rect 3396 2767 3403 2993
rect 3455 2958 3463 2982
rect 3393 2753 3407 2767
rect 3436 2727 3443 2933
rect 3496 2783 3503 3013
rect 3516 2803 3523 3233
rect 3556 3223 3563 3473
rect 3596 3327 3603 3493
rect 3636 3323 3643 3633
rect 3656 3547 3663 3573
rect 3676 3527 3683 3553
rect 3673 3513 3687 3527
rect 3696 3487 3703 3673
rect 3756 3547 3763 3713
rect 3776 3687 3783 3893
rect 3796 3687 3803 4413
rect 3816 4207 3823 4433
rect 3857 4238 3865 4262
rect 3836 4187 3843 4193
rect 3833 4173 3847 4187
rect 3857 4144 3865 4224
rect 3876 4187 3883 4453
rect 3956 4387 3963 4533
rect 3936 4183 3943 4213
rect 3953 4183 3967 4187
rect 3936 4176 3967 4183
rect 3953 4173 3967 4176
rect 3876 4087 3883 4173
rect 3916 4147 3923 4173
rect 3856 4027 3863 4033
rect 3853 4013 3867 4027
rect 3873 3973 3887 3987
rect 3936 4007 3943 4033
rect 3976 4023 3983 4513
rect 3996 4463 4003 4616
rect 4013 4463 4027 4467
rect 3996 4456 4027 4463
rect 4013 4453 4027 4456
rect 3996 4144 4004 4256
rect 4016 4167 4023 4453
rect 4036 4407 4043 4553
rect 4056 4427 4063 4573
rect 4076 4487 4083 4623
rect 4116 4587 4123 4623
rect 4136 4507 4143 4573
rect 4156 4567 4163 4623
rect 4196 4547 4203 4623
rect 4236 4587 4243 4623
rect 4256 4616 4283 4623
rect 4213 4503 4227 4507
rect 4196 4496 4227 4503
rect 4073 4473 4087 4487
rect 4096 4476 4113 4483
rect 4096 4447 4103 4476
rect 4156 4467 4163 4493
rect 4133 4433 4147 4447
rect 4153 4453 4167 4467
rect 4096 4307 4103 4433
rect 4136 4307 4143 4433
rect 4196 4407 4203 4496
rect 4213 4493 4227 4496
rect 4036 4107 4043 4293
rect 4196 4247 4203 4393
rect 4093 4173 4107 4187
rect 4136 4183 4143 4213
rect 4216 4207 4223 4233
rect 4153 4183 4167 4187
rect 4136 4176 4167 4183
rect 4213 4193 4227 4207
rect 4153 4173 4167 4176
rect 4096 4067 4103 4173
rect 4233 4173 4247 4187
rect 4196 4067 4203 4153
rect 4236 4123 4243 4173
rect 4256 4163 4263 4616
rect 4316 4587 4323 4623
rect 4556 4616 4583 4623
rect 4636 4616 4663 4623
rect 4336 4467 4343 4493
rect 4333 4453 4347 4467
rect 4256 4156 4283 4163
rect 4236 4116 4263 4123
rect 3956 4016 3983 4023
rect 3933 3993 3947 4007
rect 3856 3947 3863 3973
rect 3876 3927 3883 3973
rect 3816 3667 3823 3913
rect 3836 3664 3844 3776
rect 3896 3683 3903 3713
rect 3913 3693 3927 3707
rect 3876 3676 3903 3683
rect 3816 3527 3823 3593
rect 3773 3523 3787 3527
rect 3756 3516 3787 3523
rect 3756 3507 3763 3516
rect 3773 3513 3787 3516
rect 3813 3513 3827 3527
rect 3833 3493 3847 3507
rect 3836 3467 3843 3493
rect 3776 3327 3783 3453
rect 3636 3316 3663 3323
rect 3596 3307 3603 3313
rect 3576 3267 3583 3293
rect 3573 3253 3587 3267
rect 3536 3216 3563 3223
rect 3536 3027 3543 3216
rect 3636 3147 3643 3293
rect 3656 3267 3663 3316
rect 3776 3267 3783 3313
rect 3653 3253 3667 3267
rect 3673 3233 3687 3247
rect 3733 3263 3747 3267
rect 3716 3256 3747 3263
rect 3556 2964 3564 3076
rect 3516 2796 3543 2803
rect 3536 2787 3543 2796
rect 3496 2776 3523 2783
rect 3453 2733 3467 2747
rect 3416 2567 3423 2713
rect 3456 2687 3463 2733
rect 3473 2713 3487 2727
rect 3476 2647 3483 2713
rect 3456 2567 3463 2633
rect 3476 2567 3483 2593
rect 3496 2567 3503 2693
rect 3333 2553 3347 2567
rect 3273 2513 3287 2527
rect 3353 2533 3367 2547
rect 3373 2553 3387 2567
rect 3413 2553 3427 2567
rect 3453 2553 3467 2567
rect 3493 2553 3507 2567
rect 3276 2507 3283 2513
rect 3277 2318 3285 2342
rect 3133 2103 3147 2107
rect 3116 2096 3147 2103
rect 3133 2093 3147 2096
rect 3033 2083 3047 2087
rect 3056 2083 3063 2093
rect 3033 2076 3063 2083
rect 3033 2073 3047 2076
rect 3015 1998 3023 2022
rect 3056 1827 3063 2076
rect 3176 2087 3183 2173
rect 3196 2107 3203 2113
rect 3193 2093 3207 2107
rect 3113 2053 3127 2067
rect 3216 2087 3223 2093
rect 3213 2073 3227 2087
rect 3116 2047 3123 2053
rect 3136 2007 3143 2053
rect 3117 1838 3125 1862
rect 3013 1773 3027 1787
rect 3016 1627 3023 1773
rect 3076 1627 3083 1773
rect 3117 1744 3125 1824
rect 3136 1707 3143 1813
rect 3156 1783 3163 1853
rect 3173 1783 3187 1787
rect 3156 1776 3187 1783
rect 3173 1773 3187 1776
rect 3213 1773 3227 1787
rect 3216 1647 3223 1773
rect 3013 1623 3027 1627
rect 3013 1616 3043 1623
rect 3013 1613 3027 1616
rect 3036 1423 3043 1616
rect 3073 1613 3087 1627
rect 3136 1607 3143 1633
rect 3236 1607 3243 2253
rect 3277 2224 3285 2304
rect 3296 2207 3303 2313
rect 3333 2253 3347 2267
rect 3336 2247 3343 2253
rect 3356 2227 3363 2533
rect 3396 2527 3403 2533
rect 3416 2224 3424 2336
rect 3256 2067 3263 2153
rect 3276 2087 3283 2133
rect 3273 2073 3287 2087
rect 3353 2083 3367 2087
rect 3353 2076 3383 2083
rect 3353 2073 3367 2076
rect 3256 1744 3264 1856
rect 3133 1593 3147 1607
rect 3176 1547 3183 1593
rect 3193 1553 3207 1567
rect 3196 1547 3203 1553
rect 3016 1416 3043 1423
rect 2933 1293 2947 1307
rect 2973 1293 2987 1307
rect 2936 1267 2943 1293
rect 2976 1287 2983 1293
rect 2976 1167 2983 1273
rect 2955 1076 2963 1156
rect 2996 1147 3003 1313
rect 2996 1083 3003 1133
rect 3016 1127 3023 1416
rect 3256 1387 3263 1693
rect 3035 1358 3043 1382
rect 3035 1264 3043 1344
rect 3013 1083 3027 1087
rect 2996 1076 3027 1083
rect 3053 1083 3067 1087
rect 3076 1083 3083 1293
rect 3096 1283 3103 1333
rect 3153 1303 3167 1307
rect 3176 1303 3183 1353
rect 3216 1327 3223 1333
rect 3256 1327 3263 1353
rect 3153 1296 3183 1303
rect 3153 1293 3167 1296
rect 3193 1293 3207 1307
rect 3213 1313 3227 1327
rect 3253 1313 3267 1327
rect 3133 1283 3147 1287
rect 3096 1276 3147 1283
rect 3133 1273 3147 1276
rect 3196 1267 3203 1293
rect 3233 1273 3247 1287
rect 3236 1267 3243 1273
rect 3276 1207 3283 1933
rect 3336 1847 3343 2053
rect 3376 2047 3383 2076
rect 3416 2004 3424 2116
rect 3436 2027 3443 2513
rect 3296 1783 3303 1833
rect 3456 1827 3463 1833
rect 3313 1783 3327 1787
rect 3296 1776 3327 1783
rect 3453 1813 3467 1827
rect 3313 1773 3327 1776
rect 3353 1773 3367 1787
rect 3356 1747 3363 1773
rect 3316 1587 3323 1633
rect 3336 1607 3343 1653
rect 3293 1553 3307 1567
rect 3313 1573 3327 1587
rect 3296 1527 3303 1553
rect 3336 1547 3343 1553
rect 3136 1127 3143 1153
rect 3176 1127 3183 1133
rect 3216 1127 3223 1133
rect 3133 1113 3147 1127
rect 3013 1073 3027 1076
rect 3053 1076 3083 1083
rect 3153 1093 3167 1107
rect 3173 1113 3187 1127
rect 3213 1113 3227 1127
rect 3156 1083 3163 1093
rect 3156 1076 3183 1083
rect 3053 1073 3067 1076
rect 2955 1038 2963 1062
rect 2593 853 2607 867
rect 2596 847 2603 853
rect 2613 833 2627 847
rect 2576 807 2583 833
rect 2596 763 2603 833
rect 2616 827 2623 833
rect 2616 783 2623 813
rect 2896 847 2903 853
rect 2873 813 2887 827
rect 2893 833 2907 847
rect 2616 776 2643 783
rect 2596 756 2623 763
rect 2456 627 2463 653
rect 2476 627 2483 633
rect 2536 627 2543 713
rect 2576 627 2583 733
rect 2433 613 2447 627
rect 2533 613 2547 627
rect 2336 387 2343 393
rect 2293 383 2307 387
rect 2276 376 2307 383
rect 2213 333 2227 347
rect 2276 347 2283 376
rect 2293 373 2307 376
rect 2313 353 2327 367
rect 2316 347 2323 353
rect 2196 287 2203 333
rect 2216 327 2223 333
rect 2253 333 2267 347
rect 2233 313 2247 327
rect 2136 167 2143 213
rect 2133 153 2147 167
rect 2156 27 2163 193
rect 2176 147 2183 193
rect 2196 147 2203 213
rect 2236 163 2243 313
rect 2256 307 2263 333
rect 2393 333 2407 347
rect 2396 307 2403 333
rect 2256 207 2263 273
rect 2256 183 2263 193
rect 2356 187 2363 193
rect 2256 176 2283 183
rect 2276 167 2283 176
rect 2356 167 2363 173
rect 2396 167 2403 253
rect 2416 207 2423 413
rect 2453 373 2467 387
rect 2436 167 2443 333
rect 2456 227 2463 373
rect 2473 353 2487 367
rect 2476 347 2483 353
rect 2516 167 2523 613
rect 2573 613 2587 627
rect 2593 603 2607 607
rect 2616 603 2623 756
rect 2593 596 2623 603
rect 2593 593 2607 596
rect 2636 427 2643 776
rect 2696 627 2703 633
rect 2653 613 2667 627
rect 2693 613 2707 627
rect 2656 607 2663 613
rect 2676 547 2683 613
rect 2753 593 2767 607
rect 2536 307 2543 373
rect 2556 367 2563 413
rect 2576 367 2583 393
rect 2613 383 2627 387
rect 2596 376 2627 383
rect 2553 353 2567 367
rect 2573 323 2587 327
rect 2596 323 2603 376
rect 2613 373 2627 376
rect 2653 373 2667 387
rect 2573 316 2603 323
rect 2573 313 2587 316
rect 2556 187 2563 193
rect 2553 173 2567 187
rect 2236 156 2263 163
rect 2216 147 2223 153
rect 2213 133 2227 147
rect 2196 127 2203 133
rect 2193 113 2207 127
rect 2256 127 2263 156
rect 2273 153 2287 167
rect 2293 133 2307 147
rect 2353 153 2367 167
rect 2393 153 2407 167
rect 2433 153 2447 167
rect 2513 153 2527 167
rect 2453 143 2467 147
rect 2453 136 2483 143
rect 2596 167 2603 173
rect 2636 167 2643 353
rect 2656 327 2663 373
rect 2696 367 2703 393
rect 2736 387 2743 533
rect 2756 407 2763 593
rect 2736 367 2743 373
rect 2776 367 2783 633
rect 2836 564 2844 676
rect 2876 647 2883 813
rect 2916 647 2923 713
rect 2936 647 2943 853
rect 2996 767 3003 1053
rect 3176 847 3183 1076
rect 3013 813 3027 827
rect 3173 843 3187 847
rect 3016 807 3023 813
rect 3033 793 3047 807
rect 2873 633 2887 647
rect 2913 633 2927 647
rect 2693 353 2707 367
rect 2733 353 2747 367
rect 2856 327 2863 373
rect 2876 347 2883 413
rect 2936 387 2943 633
rect 2453 133 2467 136
rect 2233 113 2247 127
rect 2236 107 2243 113
rect 2296 87 2303 133
rect 2476 107 2483 136
rect 2533 133 2547 147
rect 2613 133 2627 147
rect 2633 153 2647 167
rect 2656 147 2663 253
rect 2696 187 2703 253
rect 2716 243 2723 313
rect 2956 247 2963 713
rect 2975 596 2983 676
rect 2993 643 3007 647
rect 3016 643 3023 793
rect 3036 667 3043 793
rect 3076 787 3083 833
rect 3093 813 3107 827
rect 3096 807 3103 813
rect 3133 813 3147 827
rect 3173 836 3203 843
rect 3173 833 3187 836
rect 3113 793 3127 807
rect 3116 787 3123 793
rect 3136 787 3143 813
rect 3196 787 3203 836
rect 3213 813 3227 827
rect 3273 833 3287 847
rect 3036 647 3043 653
rect 3076 647 3083 753
rect 3116 663 3123 773
rect 3216 667 3223 813
rect 3276 667 3283 833
rect 3133 663 3147 667
rect 3116 656 3147 663
rect 3133 653 3147 656
rect 2993 636 3023 643
rect 2993 633 3007 636
rect 3033 633 3047 647
rect 3053 613 3067 627
rect 3073 633 3087 647
rect 3056 607 3063 613
rect 2975 558 2983 582
rect 3016 367 3023 373
rect 2973 353 2987 367
rect 2976 307 2983 353
rect 2993 333 3007 347
rect 3013 353 3027 367
rect 3033 333 3047 347
rect 2716 236 2743 243
rect 2693 173 2707 187
rect 2653 133 2667 147
rect 2536 127 2543 133
rect 2616 127 2623 133
rect 2736 87 2743 236
rect 2776 167 2783 193
rect 2776 127 2783 153
rect 2773 113 2787 127
rect 2813 113 2827 127
rect 2816 87 2823 113
rect 2956 84 2964 196
rect 2996 167 3003 333
rect 3016 183 3023 233
rect 3036 207 3043 333
rect 3056 327 3063 593
rect 3176 587 3183 633
rect 3213 613 3227 627
rect 3216 587 3223 613
rect 3236 607 3243 653
rect 3296 647 3303 1373
rect 3316 1264 3324 1376
rect 3336 1147 3343 1533
rect 3356 1527 3363 1613
rect 3376 1607 3383 1773
rect 3396 1607 3403 1613
rect 3393 1593 3407 1607
rect 3413 1573 3427 1587
rect 3416 1567 3423 1573
rect 3353 1293 3367 1307
rect 3356 1247 3363 1293
rect 3376 1223 3383 1513
rect 3456 1507 3463 1753
rect 3476 1727 3483 2553
rect 3516 2527 3523 2776
rect 3556 2767 3563 2773
rect 3533 2733 3547 2747
rect 3553 2753 3567 2767
rect 3536 2667 3543 2733
rect 3536 2367 3543 2613
rect 3553 2563 3567 2567
rect 3576 2563 3583 3133
rect 3636 3047 3643 3093
rect 3676 3067 3683 3233
rect 3716 3107 3723 3256
rect 3733 3253 3747 3256
rect 3753 3233 3767 3247
rect 3773 3253 3787 3267
rect 3756 3227 3763 3233
rect 3813 3213 3827 3227
rect 3836 3223 3843 3433
rect 3876 3407 3883 3676
rect 3916 3587 3923 3693
rect 3956 3547 3963 4016
rect 3976 3996 3993 4003
rect 3976 3967 3983 3996
rect 4036 4007 4043 4053
rect 4033 3993 4047 4007
rect 4076 3963 4083 4053
rect 4096 4047 4103 4053
rect 4093 3963 4107 3967
rect 4136 3963 4143 4053
rect 4156 4007 4163 4013
rect 4153 3993 4167 4007
rect 4216 3987 4223 4093
rect 4076 3956 4107 3963
rect 4093 3953 4107 3956
rect 4116 3956 4143 3963
rect 3975 3758 3983 3782
rect 3975 3664 3983 3744
rect 3993 3703 4007 3707
rect 3993 3696 4023 3703
rect 3993 3693 4007 3696
rect 3916 3507 3923 3533
rect 3973 3513 3987 3527
rect 3893 3473 3907 3487
rect 3913 3493 3927 3507
rect 3933 3473 3947 3487
rect 3896 3467 3903 3473
rect 3936 3467 3943 3473
rect 3956 3287 3963 3513
rect 3976 3287 3983 3513
rect 3997 3476 4005 3556
rect 4016 3467 4023 3696
rect 4033 3693 4047 3707
rect 4056 3703 4063 3833
rect 4073 3703 4087 3707
rect 4056 3696 4087 3703
rect 4073 3693 4087 3696
rect 4116 3703 4123 3956
rect 4236 3867 4243 4093
rect 4256 3747 4263 4116
rect 4276 4087 4283 4156
rect 4296 4107 4303 4433
rect 4356 4227 4363 4573
rect 4393 4473 4407 4487
rect 4396 4407 4403 4473
rect 4417 4436 4425 4516
rect 4473 4483 4487 4487
rect 4473 4476 4503 4483
rect 4473 4473 4487 4476
rect 4417 4398 4425 4422
rect 4316 4143 4323 4193
rect 4333 4173 4347 4187
rect 4336 4167 4343 4173
rect 4413 4173 4427 4187
rect 4353 4153 4367 4167
rect 4356 4143 4363 4153
rect 4316 4136 4363 4143
rect 4376 4127 4383 4173
rect 4416 4127 4423 4173
rect 4496 4147 4503 4476
rect 4556 4404 4564 4516
rect 4537 4238 4545 4262
rect 4537 4144 4545 4224
rect 4336 4027 4343 4073
rect 4393 4023 4407 4027
rect 4393 4016 4423 4023
rect 4393 4013 4407 4016
rect 4333 4003 4347 4007
rect 4276 3987 4283 3993
rect 4273 3973 4287 3987
rect 4333 3996 4363 4003
rect 4333 3993 4347 3996
rect 4356 3983 4363 3996
rect 4416 4003 4423 4016
rect 4433 4003 4447 4007
rect 4416 3996 4447 4003
rect 4433 3993 4447 3996
rect 4373 3983 4387 3987
rect 4356 3976 4387 3983
rect 4373 3973 4387 3976
rect 4133 3703 4147 3707
rect 4116 3696 4147 3703
rect 4036 3567 4043 3693
rect 3997 3438 4005 3462
rect 3853 3223 3867 3227
rect 3836 3216 3867 3223
rect 3853 3213 3867 3216
rect 3816 3167 3823 3213
rect 3716 3087 3723 3093
rect 3593 3043 3607 3047
rect 3593 3036 3623 3043
rect 3593 3033 3607 3036
rect 3616 3027 3623 3036
rect 3596 2747 3603 2773
rect 3616 2704 3624 2816
rect 3553 2556 3583 2563
rect 3553 2553 3567 2556
rect 3576 2507 3583 2556
rect 3536 2287 3543 2353
rect 3556 2307 3563 2493
rect 3533 2273 3547 2287
rect 3553 2263 3567 2267
rect 3576 2263 3583 2353
rect 3616 2287 3623 2633
rect 3636 2327 3643 2873
rect 3656 2787 3663 2993
rect 3676 2867 3683 3033
rect 3695 2996 3703 3076
rect 3776 3067 3783 3073
rect 3773 3053 3787 3067
rect 3716 3007 3723 3033
rect 3695 2958 3703 2982
rect 3676 2743 3683 2853
rect 3693 2743 3707 2747
rect 3676 2736 3707 2743
rect 3693 2733 3707 2736
rect 3656 2484 3664 2596
rect 3676 2367 3683 2593
rect 3656 2287 3663 2313
rect 3553 2256 3583 2263
rect 3553 2253 3567 2256
rect 3496 2087 3503 2233
rect 3493 2073 3507 2087
rect 3496 1767 3503 2013
rect 3516 1827 3523 2213
rect 3576 2187 3583 2256
rect 3596 2247 3603 2253
rect 3613 2233 3627 2247
rect 3536 2087 3543 2113
rect 3555 2036 3563 2116
rect 3555 1998 3563 2022
rect 3537 1838 3545 1862
rect 3516 1787 3523 1813
rect 3513 1773 3527 1787
rect 3537 1744 3545 1824
rect 3476 1547 3483 1593
rect 3496 1524 3504 1636
rect 3393 1293 3407 1307
rect 3396 1287 3403 1293
rect 3396 1247 3403 1273
rect 3356 1216 3383 1223
rect 3336 1127 3343 1133
rect 3333 1113 3347 1127
rect 3356 1083 3363 1216
rect 3376 1187 3383 1193
rect 3376 1127 3383 1173
rect 3373 1123 3387 1127
rect 3393 1123 3407 1127
rect 3373 1116 3407 1123
rect 3373 1113 3387 1116
rect 3393 1113 3407 1116
rect 3416 1107 3423 1493
rect 3455 1358 3463 1382
rect 3455 1264 3463 1344
rect 3433 1123 3447 1127
rect 3456 1123 3463 1213
rect 3433 1116 3463 1123
rect 3433 1113 3447 1116
rect 3356 1076 3383 1083
rect 3376 847 3383 1076
rect 3437 878 3445 902
rect 3396 767 3403 853
rect 3437 784 3445 864
rect 3256 627 3263 633
rect 3253 613 3267 627
rect 3276 607 3283 613
rect 3273 593 3287 607
rect 3313 603 3327 607
rect 3336 603 3343 753
rect 3313 596 3343 603
rect 3313 593 3327 596
rect 3356 387 3363 673
rect 3456 667 3463 1116
rect 3476 827 3483 1153
rect 3493 813 3507 827
rect 3496 807 3503 813
rect 3496 727 3503 793
rect 3516 687 3523 1633
rect 3536 1607 3543 1613
rect 3533 1593 3547 1607
rect 3556 1603 3563 1853
rect 3596 1823 3603 2193
rect 3616 2107 3623 2233
rect 3633 2053 3647 2067
rect 3676 2067 3683 2133
rect 3673 2053 3687 2067
rect 3636 2007 3643 2053
rect 3576 1816 3603 1823
rect 3576 1783 3583 1816
rect 3593 1783 3607 1787
rect 3576 1776 3607 1783
rect 3593 1773 3607 1776
rect 3616 1763 3623 1933
rect 3633 1773 3647 1787
rect 3596 1756 3623 1763
rect 3576 1727 3583 1753
rect 3576 1627 3583 1713
rect 3573 1603 3587 1607
rect 3556 1596 3587 1603
rect 3573 1593 3587 1596
rect 3576 1127 3583 1553
rect 3596 1467 3603 1756
rect 3636 1747 3643 1773
rect 3616 1507 3623 1673
rect 3656 1647 3663 1853
rect 3676 1744 3684 1856
rect 3635 1556 3643 1636
rect 3696 1627 3703 2353
rect 3716 2327 3723 2973
rect 3776 2927 3783 3013
rect 3816 2967 3823 3013
rect 3736 2707 3743 2913
rect 3836 2887 3843 3153
rect 3856 3047 3863 3113
rect 3876 3047 3883 3253
rect 3896 3067 3903 3273
rect 3916 3267 3923 3273
rect 3913 3253 3927 3267
rect 3953 3263 3967 3267
rect 3933 3233 3947 3247
rect 3953 3256 3983 3263
rect 3953 3253 3967 3256
rect 3916 3047 3923 3133
rect 3873 3033 3887 3047
rect 3913 3033 3927 3047
rect 3936 3023 3943 3233
rect 3956 3047 3963 3213
rect 3976 3187 3983 3256
rect 4016 3247 4023 3273
rect 4036 3267 4043 3533
rect 4056 3527 4063 3573
rect 4076 3447 4083 3673
rect 4116 3667 4123 3696
rect 4133 3693 4147 3696
rect 4173 3693 4187 3707
rect 4153 3673 4167 3687
rect 4096 3527 4103 3593
rect 4093 3513 4107 3527
rect 3976 3087 3983 3173
rect 3996 3147 4003 3213
rect 4033 3213 4047 3227
rect 4053 3213 4067 3227
rect 4016 3127 4023 3153
rect 3996 3063 4003 3113
rect 4036 3087 4043 3213
rect 4056 3167 4063 3213
rect 4076 3127 4083 3313
rect 4116 3207 4123 3653
rect 4156 3627 4163 3673
rect 4176 3647 4183 3693
rect 4213 3673 4227 3687
rect 4136 3444 4144 3556
rect 4156 3427 4163 3553
rect 4176 3247 4183 3593
rect 4153 3243 4167 3247
rect 4136 3236 4167 3243
rect 3976 3056 4003 3063
rect 3976 3047 3983 3056
rect 4016 3047 4023 3073
rect 4036 3047 4043 3073
rect 3973 3033 3987 3047
rect 3953 3023 3967 3027
rect 3936 3016 3967 3023
rect 3953 3013 3967 3016
rect 4013 3033 4027 3047
rect 4033 3033 4047 3047
rect 4096 3027 4103 3053
rect 4116 3027 4123 3093
rect 4136 3087 4143 3236
rect 4153 3233 4167 3236
rect 4196 3227 4203 3673
rect 4216 3667 4223 3673
rect 4276 3627 4283 3713
rect 4296 3703 4303 3853
rect 4316 3847 4323 3973
rect 4337 3758 4345 3782
rect 4313 3703 4327 3707
rect 4296 3696 4327 3703
rect 4296 3647 4303 3696
rect 4313 3693 4327 3696
rect 4337 3664 4345 3744
rect 4213 3513 4227 3527
rect 4216 3427 4223 3513
rect 4237 3476 4245 3556
rect 4237 3438 4245 3462
rect 4316 3267 4323 3613
rect 4356 3607 4363 3953
rect 4376 3607 4383 3973
rect 4393 3693 4407 3707
rect 4333 3523 4347 3527
rect 4333 3516 4363 3523
rect 4333 3513 4347 3516
rect 4356 3467 4363 3516
rect 4336 3267 4343 3453
rect 4376 3444 4384 3556
rect 4396 3527 4403 3693
rect 4416 3627 4423 3973
rect 4457 3956 4465 4036
rect 4516 4007 4523 4133
rect 4556 4103 4563 4233
rect 4536 4096 4563 4103
rect 4513 3993 4527 4007
rect 4457 3918 4465 3942
rect 4476 3664 4484 3776
rect 4536 3767 4543 4096
rect 4576 3963 4583 4616
rect 4616 4487 4623 4513
rect 4656 4487 4663 4616
rect 4613 4473 4627 4487
rect 4653 4473 4667 4487
rect 4593 4173 4607 4187
rect 4596 4147 4603 4173
rect 4556 3956 4583 3963
rect 4396 3507 4403 3513
rect 4416 3287 4423 3593
rect 4456 3307 4463 3493
rect 4476 3283 4483 3513
rect 4496 3327 4503 3753
rect 4533 3693 4547 3707
rect 4556 3703 4563 3956
rect 4596 3924 4604 4036
rect 4573 3703 4587 3707
rect 4556 3696 4587 3703
rect 4573 3693 4587 3696
rect 4456 3276 4483 3283
rect 4213 3233 4227 3247
rect 4173 3193 4187 3207
rect 4216 3203 4223 3233
rect 4313 3243 4327 3247
rect 4296 3236 4327 3243
rect 4216 3196 4243 3203
rect 4176 3187 4183 3193
rect 4136 3047 4143 3073
rect 4133 3033 4147 3047
rect 4093 3013 4107 3027
rect 4153 3013 4167 3027
rect 4196 3027 4203 3053
rect 4193 3013 4207 3027
rect 3755 2798 3763 2822
rect 3755 2704 3763 2784
rect 3776 2747 3783 2813
rect 3773 2733 3787 2747
rect 3796 2667 3803 2773
rect 3733 2563 3747 2567
rect 3733 2556 3763 2563
rect 3733 2553 3747 2556
rect 3716 1947 3723 2233
rect 3736 1823 3743 2273
rect 3756 2207 3763 2556
rect 3776 2547 3783 2613
rect 3816 2607 3823 2833
rect 3856 2767 3863 2793
rect 3896 2767 3903 2773
rect 3833 2733 3847 2747
rect 3853 2753 3867 2767
rect 3893 2753 3907 2767
rect 3913 2733 3927 2747
rect 3836 2727 3843 2733
rect 3916 2723 3923 2733
rect 3896 2716 3923 2723
rect 3795 2516 3803 2596
rect 3813 2553 3827 2567
rect 3816 2507 3823 2553
rect 3795 2478 3803 2502
rect 3776 2327 3783 2393
rect 3816 2307 3823 2373
rect 3793 2273 3807 2287
rect 3756 2004 3764 2116
rect 3776 1823 3783 2253
rect 3796 2147 3803 2273
rect 3836 2263 3843 2713
rect 3896 2707 3903 2716
rect 3936 2707 3943 2813
rect 3976 2767 3983 2993
rect 4036 2767 4043 2813
rect 3953 2733 3967 2747
rect 3856 2487 3863 2693
rect 3916 2587 3923 2593
rect 3956 2587 3963 2733
rect 3993 2733 4007 2747
rect 4013 2733 4027 2747
rect 4033 2753 4047 2767
rect 4073 2753 4087 2767
rect 3996 2707 4003 2733
rect 4016 2727 4023 2733
rect 3996 2647 4003 2693
rect 4056 2627 4063 2713
rect 4076 2707 4083 2753
rect 3976 2587 3983 2613
rect 4096 2607 4103 2973
rect 4116 2727 4123 2993
rect 4136 2827 4143 2993
rect 4156 2967 4163 3013
rect 4176 2767 4183 2993
rect 4216 2787 4223 3153
rect 4236 3127 4243 3196
rect 4256 3167 4263 3193
rect 4256 3063 4263 3133
rect 4276 3087 4283 3193
rect 4296 3147 4303 3236
rect 4313 3233 4327 3236
rect 4353 3213 4367 3227
rect 4393 3213 4407 3227
rect 4256 3056 4283 3063
rect 4253 3023 4267 3027
rect 4276 3023 4283 3056
rect 4296 3047 4303 3113
rect 4336 3083 4343 3193
rect 4356 3187 4363 3213
rect 4356 3127 4363 3173
rect 4396 3167 4403 3213
rect 4336 3076 4363 3083
rect 4253 3016 4283 3023
rect 4253 3013 4267 3016
rect 4236 2947 4243 3013
rect 4256 2996 4273 3003
rect 4256 2847 4263 2996
rect 4316 3007 4323 3073
rect 4336 3027 4343 3053
rect 4356 3047 4363 3076
rect 4333 3013 4347 3027
rect 4313 2993 4327 3007
rect 4276 2927 4283 2973
rect 4153 2733 4167 2747
rect 4173 2753 4187 2767
rect 4193 2733 4207 2747
rect 4213 2733 4227 2747
rect 3913 2573 3927 2587
rect 3973 2573 3987 2587
rect 3936 2487 3943 2533
rect 3876 2287 3883 2353
rect 3936 2307 3943 2473
rect 3956 2307 3963 2473
rect 3976 2327 3983 2533
rect 4016 2407 4023 2593
rect 4036 2507 4043 2553
rect 4053 2533 4067 2547
rect 4056 2527 4063 2533
rect 4076 2467 4083 2573
rect 3996 2287 4003 2373
rect 4056 2307 4063 2433
rect 3853 2263 3867 2267
rect 3836 2256 3867 2263
rect 3873 2273 3887 2287
rect 3853 2253 3867 2256
rect 3893 2253 3907 2267
rect 3816 2147 3823 2253
rect 3856 2247 3863 2253
rect 3896 2243 3903 2253
rect 3896 2236 3933 2243
rect 3836 2107 3843 2193
rect 3816 2027 3823 2093
rect 3836 2087 3843 2093
rect 3833 2073 3847 2087
rect 3716 1816 3743 1823
rect 3756 1816 3783 1823
rect 3693 1623 3707 1627
rect 3653 1603 3667 1607
rect 3676 1616 3707 1623
rect 3716 1623 3723 1816
rect 3733 1773 3747 1787
rect 3736 1767 3743 1773
rect 3756 1767 3763 1816
rect 3796 1743 3803 2013
rect 3816 1823 3823 1833
rect 3876 1827 3883 2073
rect 3895 2036 3903 2116
rect 3913 2083 3927 2087
rect 3936 2083 3943 2133
rect 3913 2076 3943 2083
rect 3913 2073 3927 2076
rect 3895 1998 3903 2022
rect 3833 1823 3847 1827
rect 3816 1816 3847 1823
rect 3816 1787 3823 1816
rect 3833 1813 3847 1816
rect 3873 1813 3887 1827
rect 3776 1736 3803 1743
rect 3776 1647 3783 1736
rect 3796 1687 3803 1713
rect 3796 1627 3803 1673
rect 3716 1616 3743 1623
rect 3676 1603 3683 1616
rect 3653 1596 3683 1603
rect 3693 1613 3707 1616
rect 3653 1593 3667 1596
rect 3713 1573 3727 1587
rect 3716 1547 3723 1573
rect 3635 1518 3643 1542
rect 3616 1327 3623 1493
rect 3596 1263 3603 1273
rect 3636 1263 3643 1273
rect 3596 1256 3643 1263
rect 3576 784 3584 896
rect 3596 827 3603 1113
rect 3616 1103 3623 1233
rect 3633 1103 3647 1107
rect 3616 1096 3647 1103
rect 3633 1093 3647 1096
rect 3636 867 3643 1093
rect 3656 987 3663 1453
rect 3736 1347 3743 1616
rect 3793 1613 3807 1627
rect 3756 1583 3763 1613
rect 3773 1583 3787 1587
rect 3756 1576 3787 1583
rect 3773 1573 3787 1576
rect 3673 1293 3687 1307
rect 3676 1287 3683 1293
rect 3716 1283 3723 1293
rect 3733 1283 3747 1287
rect 3716 1276 3747 1283
rect 3733 1273 3747 1276
rect 3673 813 3687 827
rect 3676 687 3683 813
rect 3716 807 3723 853
rect 3416 603 3423 633
rect 3433 603 3447 607
rect 3416 596 3447 603
rect 3473 603 3487 607
rect 3496 603 3503 653
rect 3576 647 3583 653
rect 3433 593 3447 596
rect 3473 596 3503 603
rect 3573 633 3587 647
rect 3473 593 3487 596
rect 3476 427 3483 593
rect 3636 564 3644 676
rect 3716 647 3723 793
rect 3756 784 3764 896
rect 3776 727 3783 1553
rect 3796 1287 3803 1573
rect 3816 1567 3823 1753
rect 3876 1747 3883 1773
rect 3836 1607 3843 1653
rect 3856 1607 3863 1693
rect 3896 1687 3903 1933
rect 3916 1867 3923 2053
rect 3956 1827 3963 2273
rect 3973 2253 3987 2267
rect 3993 2273 4007 2287
rect 4053 2253 4067 2267
rect 3976 2247 3983 2253
rect 4056 2243 4063 2253
rect 4007 2236 4063 2243
rect 3997 2036 4005 2116
rect 3997 1998 4005 2022
rect 3933 1783 3947 1787
rect 3927 1776 3947 1783
rect 3933 1773 3947 1776
rect 3996 1763 4003 1953
rect 4016 1947 4023 2213
rect 4036 2087 4043 2213
rect 4056 2087 4063 2093
rect 4053 2073 4067 2087
rect 4056 1807 4063 2013
rect 4076 1967 4083 2453
rect 4096 2103 4103 2493
rect 4116 2447 4123 2693
rect 4156 2687 4163 2733
rect 4196 2727 4203 2733
rect 4136 2347 4143 2653
rect 4116 2224 4124 2336
rect 4156 2303 4163 2613
rect 4136 2296 4163 2303
rect 4136 2163 4143 2296
rect 4153 2253 4167 2267
rect 4156 2247 4163 2253
rect 4136 2156 4163 2163
rect 4096 2096 4123 2103
rect 4116 1867 4123 2096
rect 4136 2004 4144 2116
rect 4156 1963 4163 2156
rect 4136 1956 4163 1963
rect 4013 1793 4027 1807
rect 3976 1756 4003 1763
rect 3896 1607 3903 1653
rect 3853 1593 3867 1607
rect 3893 1603 3907 1607
rect 3913 1603 3927 1607
rect 3893 1596 3927 1603
rect 3956 1607 3963 1713
rect 3893 1593 3907 1596
rect 3913 1593 3927 1596
rect 3953 1593 3967 1607
rect 3976 1563 3983 1756
rect 3996 1703 4003 1733
rect 4016 1727 4023 1793
rect 4053 1793 4067 1807
rect 4073 1773 4087 1787
rect 3996 1696 4023 1703
rect 4016 1627 4023 1696
rect 4013 1613 4027 1627
rect 4036 1607 4043 1753
rect 4056 1667 4063 1753
rect 4076 1747 4083 1773
rect 4093 1753 4107 1767
rect 4096 1707 4103 1753
rect 4076 1643 4083 1693
rect 4116 1667 4123 1773
rect 4056 1636 4083 1643
rect 4033 1593 4047 1607
rect 3956 1556 3983 1563
rect 3837 1358 3845 1382
rect 3956 1347 3963 1556
rect 3837 1264 3845 1344
rect 3856 1147 3863 1333
rect 3876 1267 3883 1333
rect 3893 1293 3907 1307
rect 3896 1147 3903 1293
rect 3976 1264 3984 1376
rect 4016 1207 4023 1573
rect 4056 1547 4063 1636
rect 4096 1627 4103 1653
rect 4136 1623 4143 1956
rect 4156 1807 4163 1933
rect 4153 1793 4167 1807
rect 4156 1627 4163 1653
rect 4176 1627 4183 2713
rect 4216 2647 4223 2733
rect 4253 2733 4267 2747
rect 4216 2267 4223 2533
rect 4236 2487 4243 2693
rect 4256 2527 4263 2733
rect 4276 2727 4283 2853
rect 4276 2484 4284 2596
rect 4255 2318 4263 2342
rect 4193 2263 4207 2267
rect 4193 2256 4213 2263
rect 4193 2253 4207 2256
rect 4196 2107 4203 2253
rect 4236 2183 4243 2233
rect 4255 2224 4263 2304
rect 4273 2263 4287 2267
rect 4296 2263 4303 2973
rect 4316 2707 4323 2933
rect 4336 2704 4344 2816
rect 4376 2783 4383 3133
rect 4396 3067 4403 3113
rect 4416 3087 4423 3213
rect 4436 3187 4443 3273
rect 4356 2776 4383 2783
rect 4356 2583 4363 2776
rect 4396 2647 4403 3053
rect 4416 2967 4423 3013
rect 4437 2996 4445 3076
rect 4437 2958 4445 2982
rect 4413 2733 4427 2747
rect 4416 2727 4423 2733
rect 4436 2727 4443 2873
rect 4356 2576 4383 2583
rect 4353 2563 4367 2567
rect 4336 2556 4367 2563
rect 4336 2547 4343 2556
rect 4353 2553 4367 2556
rect 4273 2256 4303 2263
rect 4273 2253 4287 2256
rect 4316 2223 4323 2513
rect 4357 2318 4365 2342
rect 4336 2267 4343 2293
rect 4333 2253 4347 2267
rect 4357 2224 4365 2304
rect 4316 2216 4343 2223
rect 4236 2176 4263 2183
rect 4256 2087 4263 2176
rect 4296 2087 4303 2133
rect 4316 2107 4323 2113
rect 4336 2107 4343 2216
rect 4376 2147 4383 2576
rect 4415 2516 4423 2596
rect 4433 2553 4447 2567
rect 4436 2547 4443 2553
rect 4415 2478 4423 2502
rect 4416 2147 4423 2253
rect 4313 2093 4327 2107
rect 4213 2083 4227 2087
rect 4196 2076 4227 2083
rect 4196 1947 4203 2076
rect 4213 2073 4227 2076
rect 4233 2053 4247 2067
rect 4253 2073 4267 2087
rect 4273 2053 4287 2067
rect 4293 2073 4307 2087
rect 4236 1927 4243 2053
rect 4116 1616 4143 1623
rect 4033 1293 4047 1307
rect 4036 1247 4043 1293
rect 3713 633 3727 647
rect 3775 596 3783 676
rect 3816 667 3823 1133
rect 3896 1107 3903 1133
rect 3833 823 3847 827
rect 3856 823 3863 1093
rect 3895 878 3903 902
rect 3833 816 3863 823
rect 3833 813 3847 816
rect 3856 807 3863 816
rect 3895 784 3903 864
rect 3916 827 3923 973
rect 3936 963 3943 1193
rect 4053 1113 4067 1127
rect 3953 1073 3967 1087
rect 3993 1083 4007 1087
rect 4016 1083 4023 1113
rect 3993 1076 4023 1083
rect 3993 1073 4007 1076
rect 3956 987 3963 1073
rect 3936 956 3963 963
rect 3913 813 3927 827
rect 3936 787 3943 853
rect 3836 647 3843 673
rect 3793 633 3807 647
rect 3833 633 3847 647
rect 3775 558 3783 582
rect 3796 547 3803 633
rect 3853 613 3867 627
rect 3476 387 3483 413
rect 3116 367 3123 373
rect 3093 333 3107 347
rect 3113 353 3127 367
rect 3253 363 3267 367
rect 3236 356 3267 363
rect 3236 347 3243 356
rect 3253 353 3267 356
rect 3213 343 3227 347
rect 3096 307 3103 333
rect 3016 176 3033 183
rect 3036 167 3043 173
rect 3076 167 3083 213
rect 2993 153 3007 167
rect 3033 153 3047 167
rect 3095 116 3103 196
rect 3136 147 3143 333
rect 3213 336 3233 343
rect 3213 333 3227 336
rect 3193 313 3207 327
rect 3333 333 3347 347
rect 3373 343 3387 347
rect 3396 343 3403 373
rect 3373 336 3403 343
rect 3373 333 3387 336
rect 3413 333 3427 347
rect 3473 363 3487 367
rect 3473 356 3503 363
rect 3473 353 3487 356
rect 3273 313 3287 327
rect 3196 287 3203 313
rect 3276 267 3283 313
rect 3336 247 3343 333
rect 3416 327 3423 333
rect 3496 307 3503 356
rect 3156 187 3163 213
rect 3153 173 3167 187
rect 3173 143 3187 147
rect 3196 143 3203 193
rect 3253 183 3267 187
rect 3253 176 3283 183
rect 3253 173 3267 176
rect 3173 136 3203 143
rect 3276 167 3283 176
rect 3173 133 3187 136
rect 3095 78 3103 102
rect 3316 84 3324 196
rect 3356 167 3363 293
rect 3516 287 3523 333
rect 3553 333 3567 347
rect 3616 347 3623 393
rect 3636 367 3643 393
rect 3796 387 3803 393
rect 3673 383 3687 387
rect 3656 376 3687 383
rect 3713 383 3727 387
rect 3633 353 3647 367
rect 3396 167 3403 173
rect 3353 153 3367 167
rect 3393 153 3407 167
rect 3455 116 3463 196
rect 3556 187 3563 333
rect 3593 333 3607 347
rect 3596 327 3603 333
rect 3656 327 3663 376
rect 3673 373 3687 376
rect 3713 376 3743 383
rect 3713 373 3727 376
rect 3573 313 3587 327
rect 3576 307 3583 313
rect 3736 307 3743 376
rect 3793 373 3807 387
rect 3553 173 3567 187
rect 3576 167 3583 253
rect 3637 116 3645 196
rect 3696 167 3703 173
rect 3736 167 3743 233
rect 3693 153 3707 167
rect 3733 153 3747 167
rect 3455 78 3463 102
rect 3637 78 3645 102
rect 3776 84 3784 196
rect 3796 147 3803 173
rect 3816 167 3823 613
rect 3856 603 3863 613
rect 3836 596 3863 603
rect 3836 367 3843 596
rect 3916 587 3923 633
rect 3936 603 3943 673
rect 3956 647 3963 956
rect 4036 867 4043 1093
rect 4056 1087 4063 1113
rect 4077 1076 4085 1156
rect 4077 1038 4085 1062
rect 4097 878 4105 902
rect 4016 847 4023 853
rect 4013 833 4027 847
rect 4033 813 4047 827
rect 4036 687 4043 813
rect 4097 784 4105 864
rect 4116 823 4123 1616
rect 4153 1613 4167 1627
rect 4196 1607 4203 1913
rect 4276 1847 4283 2053
rect 4316 2023 4323 2053
rect 4336 2047 4343 2053
rect 4316 2016 4343 2023
rect 4336 1787 4343 2016
rect 4356 1807 4363 2093
rect 4393 2083 4407 2087
rect 4376 2076 4407 2083
rect 4436 2087 4443 2513
rect 4456 2507 4463 3276
rect 4516 3267 4523 3273
rect 4513 3253 4527 3267
rect 4476 2867 4483 3073
rect 4496 3047 4503 3073
rect 4536 3063 4543 3693
rect 4593 3493 4607 3507
rect 4516 3056 4543 3063
rect 4493 3033 4507 3047
rect 4475 2798 4483 2822
rect 4475 2704 4483 2784
rect 4496 2747 4503 2773
rect 4493 2733 4507 2747
rect 4516 2687 4523 3056
rect 4556 2987 4563 3493
rect 4596 3487 4603 3493
rect 4616 3463 4623 4433
rect 4676 4307 4683 4453
rect 4693 4433 4707 4447
rect 4633 4173 4647 4187
rect 4636 4127 4643 4173
rect 4676 4144 4684 4256
rect 4653 4023 4667 4027
rect 4636 4016 4667 4023
rect 4636 3967 4643 4016
rect 4653 4013 4667 4016
rect 4636 3727 4643 3913
rect 4696 3783 4703 4433
rect 4716 3987 4723 4193
rect 4696 3776 4723 3783
rect 4696 3727 4703 3753
rect 4693 3713 4707 3727
rect 4653 3673 4667 3687
rect 4656 3667 4663 3673
rect 4596 3456 4623 3463
rect 4576 3184 4584 3296
rect 4576 2964 4584 3076
rect 4596 3007 4603 3456
rect 4613 3213 4627 3227
rect 4636 3223 4643 3293
rect 4656 3267 4663 3453
rect 4676 3287 4683 3473
rect 4716 3343 4723 3776
rect 4696 3336 4723 3343
rect 4653 3223 4667 3227
rect 4636 3216 4667 3223
rect 4616 3047 4623 3213
rect 4636 3087 4643 3216
rect 4653 3213 4667 3216
rect 4656 3107 4663 3193
rect 4656 3063 4663 3073
rect 4676 3067 4683 3233
rect 4696 3227 4703 3336
rect 4715 3278 4723 3302
rect 4636 3056 4663 3063
rect 4636 3047 4643 3056
rect 4633 3033 4647 3047
rect 4653 3013 4667 3027
rect 4696 3043 4703 3213
rect 4715 3184 4723 3264
rect 4736 3247 4743 4293
rect 4736 3087 4743 3173
rect 4696 3036 4723 3043
rect 4616 2927 4623 3013
rect 4656 3007 4663 3013
rect 4676 2807 4683 2993
rect 4556 2767 4563 2793
rect 4533 2733 4547 2747
rect 4553 2753 4567 2767
rect 4593 2753 4607 2767
rect 4536 2727 4543 2733
rect 4596 2727 4603 2753
rect 4476 2567 4483 2573
rect 4473 2553 4487 2567
rect 4493 2533 4507 2547
rect 4536 2547 4543 2553
rect 4533 2533 4547 2547
rect 4496 2487 4503 2533
rect 4556 2527 4563 2693
rect 4616 2567 4623 2793
rect 4676 2787 4683 2793
rect 4653 2753 4667 2767
rect 4673 2773 4687 2787
rect 4596 2547 4603 2553
rect 4593 2533 4607 2547
rect 4636 2527 4643 2733
rect 4656 2727 4663 2753
rect 4676 2547 4683 2733
rect 4696 2707 4703 2973
rect 4653 2513 4667 2527
rect 4673 2533 4687 2547
rect 4576 2347 4583 2513
rect 4616 2487 4623 2513
rect 4656 2507 4663 2513
rect 4496 2224 4504 2336
rect 4656 2343 4663 2493
rect 4636 2336 4663 2343
rect 4536 2167 4543 2293
rect 4576 2287 4583 2313
rect 4553 2253 4567 2267
rect 4573 2273 4587 2287
rect 4556 2187 4563 2253
rect 4636 2183 4643 2336
rect 4696 2327 4703 2473
rect 4696 2307 4703 2313
rect 4693 2293 4707 2307
rect 4636 2176 4663 2183
rect 4476 2087 4483 2113
rect 4433 2083 4447 2087
rect 4376 2067 4383 2076
rect 4393 2073 4407 2076
rect 4433 2076 4463 2083
rect 4433 2073 4447 2076
rect 4456 1823 4463 2076
rect 4473 2073 4487 2087
rect 4477 1838 4485 1862
rect 4436 1816 4463 1823
rect 4313 1773 4327 1787
rect 4356 1783 4363 1793
rect 4373 1783 4387 1787
rect 4356 1776 4387 1783
rect 4373 1773 4387 1776
rect 4273 1753 4287 1767
rect 4216 1627 4223 1693
rect 4236 1607 4243 1733
rect 4276 1707 4283 1753
rect 4133 1573 4147 1587
rect 4173 1573 4187 1587
rect 4193 1593 4207 1607
rect 4233 1603 4247 1607
rect 4216 1596 4247 1603
rect 4276 1607 4283 1653
rect 4216 1587 4223 1596
rect 4233 1593 4247 1596
rect 4273 1593 4287 1607
rect 4136 1547 4143 1573
rect 4176 1407 4183 1573
rect 4136 1347 4143 1353
rect 4176 1347 4183 1373
rect 4133 1333 4147 1347
rect 4173 1333 4187 1347
rect 4136 1127 4143 1133
rect 4176 1127 4183 1133
rect 4133 1113 4147 1127
rect 4173 1113 4187 1127
rect 4196 1087 4203 1533
rect 4216 1507 4223 1553
rect 4256 1547 4263 1573
rect 4296 1427 4303 1673
rect 4316 1667 4323 1773
rect 4336 1763 4343 1773
rect 4336 1756 4363 1763
rect 4336 1627 4343 1693
rect 4356 1627 4363 1756
rect 4313 1573 4327 1587
rect 4316 1567 4323 1573
rect 4216 1303 4223 1353
rect 4233 1303 4247 1307
rect 4216 1296 4247 1303
rect 4233 1293 4247 1296
rect 4216 1044 4224 1156
rect 4116 816 4143 823
rect 3953 603 3967 607
rect 3936 596 3967 603
rect 3953 593 3967 596
rect 3896 367 3903 413
rect 3853 353 3867 367
rect 3856 347 3863 353
rect 3873 333 3887 347
rect 3893 353 3907 367
rect 3953 363 3967 367
rect 3913 343 3927 347
rect 3936 356 3967 363
rect 3936 343 3943 356
rect 3913 336 3943 343
rect 3953 353 3967 356
rect 3913 333 3927 336
rect 3876 287 3883 333
rect 3916 267 3923 333
rect 3973 313 3987 327
rect 3976 307 3983 313
rect 3936 167 3943 293
rect 3853 143 3867 147
rect 3876 143 3883 153
rect 3853 136 3883 143
rect 3853 133 3867 136
rect 3913 133 3927 147
rect 3933 153 3947 167
rect 3956 147 3963 213
rect 3953 133 3967 147
rect 3916 127 3923 133
rect 3976 127 3983 253
rect 3996 187 4003 533
rect 4016 367 4023 653
rect 4036 607 4043 633
rect 4057 596 4065 676
rect 4057 558 4065 582
rect 4076 367 4083 773
rect 4116 647 4123 793
rect 4113 633 4127 647
rect 4096 587 4103 633
rect 4097 398 4105 422
rect 4013 353 4027 367
rect 4097 304 4105 384
rect 4116 307 4123 333
rect 4136 327 4143 816
rect 4153 813 4167 827
rect 4193 813 4207 827
rect 4156 807 4163 813
rect 4153 343 4167 347
rect 4176 343 4183 793
rect 4196 767 4203 813
rect 4236 784 4244 896
rect 4256 827 4263 1413
rect 4296 1343 4303 1393
rect 4356 1347 4363 1553
rect 4313 1343 4327 1347
rect 4296 1336 4327 1343
rect 4273 1293 4287 1307
rect 4276 1187 4283 1293
rect 4296 1127 4303 1336
rect 4313 1333 4327 1336
rect 4353 1333 4367 1347
rect 4376 1307 4383 1513
rect 4396 1387 4403 1733
rect 4416 1667 4423 1673
rect 4436 1667 4443 1816
rect 4456 1787 4463 1793
rect 4453 1773 4467 1787
rect 4477 1744 4485 1824
rect 4496 1787 4503 2053
rect 4416 1627 4423 1653
rect 4413 1613 4427 1627
rect 4456 1567 4463 1713
rect 4476 1627 4483 1693
rect 4516 1627 4523 1833
rect 4536 1823 4543 2133
rect 4556 1847 4563 2073
rect 4577 2036 4585 2116
rect 4577 1998 4585 2022
rect 4536 1816 4563 1823
rect 4533 1783 4547 1787
rect 4556 1783 4563 1816
rect 4533 1776 4563 1783
rect 4533 1773 4547 1776
rect 4596 1747 4603 2153
rect 4636 2087 4643 2133
rect 4633 2073 4647 2087
rect 4616 1744 4624 1856
rect 4656 1827 4663 2176
rect 4676 2087 4683 2253
rect 4716 2163 4723 3036
rect 4736 3027 4743 3053
rect 4736 2267 4743 2993
rect 4756 2747 4763 3493
rect 4776 3087 4783 3713
rect 4776 2927 4783 3053
rect 4696 2156 4723 2163
rect 4673 2073 4687 2087
rect 4696 1827 4703 2156
rect 4716 2004 4724 2116
rect 4693 1813 4707 1827
rect 4656 1727 4663 1813
rect 4713 1793 4727 1807
rect 4473 1613 4487 1627
rect 4476 1367 4483 1553
rect 4476 1323 4483 1353
rect 4516 1343 4523 1593
rect 4536 1583 4543 1653
rect 4553 1583 4567 1587
rect 4536 1576 4567 1583
rect 4553 1573 4567 1576
rect 4656 1587 4663 1673
rect 4676 1627 4683 1773
rect 4716 1607 4723 1793
rect 4776 1607 4783 2333
rect 4653 1573 4667 1587
rect 4647 1516 4653 1523
rect 4676 1367 4683 1593
rect 4516 1336 4543 1343
rect 4536 1327 4543 1336
rect 4493 1323 4507 1327
rect 4453 1293 4467 1307
rect 4476 1316 4507 1323
rect 4456 1267 4463 1293
rect 4396 1127 4403 1133
rect 4313 1083 4327 1087
rect 4336 1083 4343 1113
rect 4393 1113 4407 1127
rect 4313 1076 4343 1083
rect 4436 1087 4443 1153
rect 4476 1123 4483 1316
rect 4493 1313 4507 1316
rect 4513 1293 4527 1307
rect 4573 1293 4587 1307
rect 4613 1303 4627 1307
rect 4636 1303 4643 1353
rect 4496 1127 4503 1293
rect 4516 1287 4523 1293
rect 4556 1147 4563 1293
rect 4576 1287 4583 1293
rect 4613 1296 4643 1303
rect 4613 1293 4627 1296
rect 4593 1273 4607 1287
rect 4596 1267 4603 1273
rect 4536 1136 4553 1143
rect 4536 1127 4543 1136
rect 4576 1127 4583 1153
rect 4636 1127 4643 1296
rect 4456 1116 4483 1123
rect 4313 1073 4327 1076
rect 4196 564 4204 676
rect 4216 607 4223 713
rect 4236 463 4243 613
rect 4293 593 4307 607
rect 4316 603 4323 813
rect 4336 784 4344 896
rect 4373 813 4387 827
rect 4456 827 4463 1116
rect 4533 1113 4547 1127
rect 4573 1113 4587 1127
rect 4633 1103 4647 1107
rect 4656 1103 4663 1273
rect 4696 1127 4703 1353
rect 4736 1327 4743 1333
rect 4756 1327 4763 1593
rect 4776 1367 4783 1573
rect 4733 1313 4747 1327
rect 4676 1107 4683 1113
rect 4513 1073 4527 1087
rect 4616 1096 4663 1103
rect 4516 1047 4523 1073
rect 4475 878 4483 902
rect 4413 813 4427 827
rect 4376 787 4383 813
rect 4416 807 4423 813
rect 4475 784 4483 864
rect 4496 827 4503 913
rect 4556 907 4563 1073
rect 4616 927 4623 1096
rect 4633 1093 4647 1096
rect 4673 1093 4687 1107
rect 4693 1073 4707 1087
rect 4556 847 4563 893
rect 4493 813 4507 827
rect 4533 813 4547 827
rect 4553 833 4567 847
rect 4593 843 4607 847
rect 4616 843 4623 873
rect 4656 847 4663 913
rect 4676 867 4683 1053
rect 4696 1047 4703 1073
rect 4593 836 4623 843
rect 4593 833 4607 836
rect 4573 823 4587 827
rect 4573 816 4603 823
rect 4573 813 4587 816
rect 4333 603 4347 607
rect 4316 596 4347 603
rect 4373 603 4387 607
rect 4396 603 4403 673
rect 4456 647 4463 753
rect 4496 647 4503 673
rect 4453 633 4467 647
rect 4333 593 4347 596
rect 4373 596 4403 603
rect 4473 613 4487 627
rect 4493 633 4507 647
rect 4373 593 4387 596
rect 4236 456 4263 463
rect 4153 336 4183 343
rect 4153 333 4167 336
rect 4193 333 4207 347
rect 4036 167 4043 253
rect 4093 183 4107 187
rect 4056 176 4107 183
rect 4033 153 4047 167
rect 4056 147 4063 176
rect 4093 173 4107 176
rect 4116 167 4123 293
rect 4196 287 4203 333
rect 4236 304 4244 416
rect 4256 347 4263 456
rect 4296 427 4303 593
rect 4476 527 4483 613
rect 4536 427 4543 813
rect 4556 564 4564 676
rect 4596 647 4603 816
rect 4653 833 4667 847
rect 4693 843 4707 847
rect 4716 843 4723 1313
rect 4753 1283 4767 1287
rect 4776 1283 4783 1313
rect 4753 1276 4783 1283
rect 4753 1273 4767 1276
rect 4736 887 4743 1113
rect 4756 927 4763 1133
rect 4693 836 4723 843
rect 4693 833 4707 836
rect 4673 823 4687 827
rect 4673 816 4703 823
rect 4673 813 4687 816
rect 4636 647 4643 793
rect 4676 647 4683 793
rect 4696 787 4703 816
rect 4593 633 4607 647
rect 4633 643 4647 647
rect 4616 636 4647 643
rect 4176 196 4223 203
rect 4176 187 4183 196
rect 4216 183 4223 196
rect 4216 176 4243 183
rect 4176 167 4183 173
rect 4113 153 4127 167
rect 4173 153 4187 167
rect 4236 167 4243 176
rect 4276 167 4283 393
rect 4356 387 4363 393
rect 4353 373 4367 387
rect 4376 227 4383 373
rect 4393 353 4407 367
rect 4396 347 4403 353
rect 4413 333 4427 347
rect 4453 343 4467 347
rect 4476 343 4483 413
rect 4577 398 4585 422
rect 4453 336 4483 343
rect 4553 343 4567 347
rect 4453 333 4467 336
rect 4416 307 4423 333
rect 4513 323 4527 327
rect 4536 336 4567 343
rect 4536 323 4543 336
rect 4513 316 4543 323
rect 4553 333 4567 336
rect 4513 313 4527 316
rect 4233 153 4247 167
rect 4273 153 4287 167
rect 4336 123 4343 173
rect 4376 147 4383 213
rect 4353 123 4367 127
rect 4336 116 4367 123
rect 4373 133 4387 147
rect 4393 123 4407 127
rect 4416 123 4423 173
rect 4476 167 4483 313
rect 4577 304 4585 384
rect 4616 343 4623 636
rect 4633 633 4647 636
rect 4633 343 4647 347
rect 4616 336 4647 343
rect 4633 333 4647 336
rect 4516 187 4523 193
rect 4656 183 4663 633
rect 4695 596 4703 676
rect 4695 558 4703 582
rect 4673 333 4687 347
rect 4676 307 4683 333
rect 4696 263 4703 513
rect 4716 304 4724 416
rect 4696 256 4723 263
rect 4673 183 4687 187
rect 4656 176 4687 183
rect 4673 173 4687 176
rect 4516 167 4523 173
rect 4513 153 4527 167
rect 4353 113 4367 116
rect 4393 116 4423 123
rect 4393 113 4407 116
rect 4436 107 4443 133
rect 4536 123 4543 153
rect 4553 123 4567 127
rect 4536 116 4567 123
rect 4593 123 4607 127
rect 4616 123 4623 173
rect 4716 147 4723 256
rect 4756 147 4763 893
rect 4553 113 4567 116
rect 4593 116 4623 123
rect 4593 113 4607 116
rect 4713 133 4727 147
rect 4733 113 4747 127
rect 4736 107 4743 113
rect 1976 -24 1983 13
rect 2116 -24 2123 13
<< m3contact >>
rect 1233 4553 1247 4567
rect 1533 4553 1547 4567
rect 113 4533 127 4547
rect 193 4533 207 4547
rect 893 4533 907 4547
rect 33 4513 47 4527
rect 73 4493 87 4507
rect 93 4453 107 4467
rect 93 4413 107 4427
rect 173 4493 187 4507
rect 173 4473 187 4487
rect 153 4453 167 4467
rect 493 4513 507 4527
rect 713 4513 727 4527
rect 373 4493 387 4507
rect 433 4493 447 4507
rect 553 4493 567 4507
rect 653 4493 667 4507
rect 213 4473 227 4487
rect 173 4433 187 4447
rect 233 4453 247 4467
rect 253 4453 267 4467
rect 53 4393 67 4407
rect 113 4393 127 4407
rect 153 4413 167 4427
rect 313 4453 327 4467
rect 273 4433 287 4447
rect 193 4413 207 4427
rect 133 4353 147 4367
rect 33 4233 47 4247
rect 93 4233 107 4247
rect 73 4213 87 4227
rect 173 4393 187 4407
rect 153 4213 167 4227
rect 93 4193 107 4207
rect 73 4173 87 4187
rect 133 4193 147 4207
rect 53 4133 67 4147
rect 53 4033 67 4047
rect 113 4153 127 4167
rect 73 4013 87 4027
rect 173 4113 187 4127
rect 153 4093 167 4107
rect 153 4073 167 4087
rect 33 3953 47 3967
rect 53 3893 67 3907
rect 133 3933 147 3947
rect 353 4453 367 4467
rect 393 4473 407 4487
rect 413 4453 427 4467
rect 453 4453 467 4467
rect 473 4473 487 4487
rect 493 4453 507 4467
rect 613 4473 627 4487
rect 373 4433 387 4447
rect 333 4393 347 4407
rect 513 4433 527 4447
rect 533 4433 547 4447
rect 673 4453 687 4467
rect 693 4453 707 4467
rect 613 4433 627 4447
rect 553 4353 567 4367
rect 593 4353 607 4367
rect 453 4313 467 4327
rect 353 4273 367 4287
rect 413 4273 427 4287
rect 213 4213 227 4227
rect 233 4193 247 4207
rect 253 4173 267 4187
rect 193 4053 207 4067
rect 213 4013 227 4027
rect 313 4213 327 4227
rect 293 4173 307 4187
rect 353 4173 367 4187
rect 313 4153 327 4167
rect 293 4133 307 4147
rect 393 4173 407 4187
rect 413 4193 427 4207
rect 473 4193 487 4207
rect 513 4193 527 4207
rect 493 4173 507 4187
rect 373 4113 387 4127
rect 573 4313 587 4327
rect 653 4433 667 4447
rect 633 4413 647 4427
rect 753 4473 767 4487
rect 773 4473 787 4487
rect 833 4473 847 4487
rect 853 4473 867 4487
rect 753 4453 767 4467
rect 793 4453 807 4467
rect 813 4453 827 4467
rect 853 4453 867 4467
rect 713 4413 727 4427
rect 833 4433 847 4447
rect 873 4433 887 4447
rect 813 4413 827 4427
rect 853 4413 867 4427
rect 1053 4493 1067 4507
rect 1073 4493 1087 4507
rect 1113 4493 1127 4507
rect 1133 4493 1147 4507
rect 993 4473 1007 4487
rect 933 4453 947 4467
rect 953 4433 967 4447
rect 1033 4453 1047 4467
rect 1013 4433 1027 4447
rect 693 4393 707 4407
rect 653 4373 667 4387
rect 653 4213 667 4227
rect 693 4193 707 4207
rect 553 4153 567 4167
rect 733 4373 747 4387
rect 813 4353 827 4367
rect 793 4213 807 4227
rect 773 4193 787 4207
rect 673 4153 687 4167
rect 693 4153 707 4167
rect 713 4153 727 4167
rect 753 4153 767 4167
rect 593 4133 607 4147
rect 513 4113 527 4127
rect 593 4113 607 4127
rect 433 4093 447 4107
rect 273 4073 287 4087
rect 333 4073 347 4087
rect 293 4053 307 4067
rect 373 4033 387 4047
rect 413 4033 427 4047
rect 333 4013 347 4027
rect 193 3953 207 3967
rect 253 3973 267 3987
rect 273 3973 287 3987
rect 493 4013 507 4027
rect 153 3873 167 3887
rect 173 3873 187 3887
rect 73 3733 87 3747
rect 133 3733 147 3747
rect 53 3713 67 3727
rect 73 3693 87 3707
rect 113 3713 127 3727
rect 153 3713 167 3727
rect 153 3693 167 3707
rect 53 3673 67 3687
rect 73 3653 87 3667
rect 113 3673 127 3687
rect 53 3633 67 3647
rect 93 3633 107 3647
rect 33 3613 47 3627
rect 133 3653 147 3667
rect 93 3613 107 3627
rect 113 3613 127 3627
rect 13 3473 27 3487
rect 73 3473 87 3487
rect 13 3413 27 3427
rect 13 3393 27 3407
rect 113 3593 127 3607
rect 113 3473 127 3487
rect 33 3273 47 3287
rect 13 3193 27 3207
rect 93 3433 107 3447
rect 93 3253 107 3267
rect 113 3253 127 3267
rect 93 3213 107 3227
rect 93 3193 107 3207
rect 93 3153 107 3167
rect 133 3193 147 3207
rect 173 3653 187 3667
rect 173 3533 187 3547
rect 253 3913 267 3927
rect 353 3953 367 3967
rect 213 3713 227 3727
rect 313 3893 327 3907
rect 433 3993 447 4007
rect 513 3993 527 4007
rect 553 3973 567 3987
rect 453 3933 467 3947
rect 573 3933 587 3947
rect 433 3913 447 3927
rect 533 3913 547 3927
rect 653 4053 667 4067
rect 613 3993 627 4007
rect 633 3973 647 3987
rect 673 3973 687 3987
rect 653 3933 667 3947
rect 393 3893 407 3907
rect 533 3893 547 3907
rect 593 3893 607 3907
rect 373 3873 387 3887
rect 413 3753 427 3767
rect 393 3733 407 3747
rect 293 3713 307 3727
rect 333 3713 347 3727
rect 353 3713 367 3727
rect 353 3693 367 3707
rect 233 3673 247 3687
rect 253 3673 267 3687
rect 313 3673 327 3687
rect 233 3633 247 3647
rect 173 3233 187 3247
rect 173 3213 187 3227
rect 133 3173 147 3187
rect 153 3173 167 3187
rect 133 3133 147 3147
rect 213 3213 227 3227
rect 313 3633 327 3647
rect 293 3433 307 3447
rect 293 3393 307 3407
rect 253 3353 267 3367
rect 253 3333 267 3347
rect 233 3193 247 3207
rect 33 3033 47 3047
rect 93 3013 107 3027
rect 113 3033 127 3047
rect 33 2993 47 3007
rect 13 2933 27 2947
rect 13 2773 27 2787
rect 73 2993 87 3007
rect 153 3053 167 3067
rect 53 2973 67 2987
rect 53 2913 67 2927
rect 93 2973 107 2987
rect 73 2833 87 2847
rect 33 2753 47 2767
rect 53 2753 67 2767
rect 33 2713 47 2727
rect 13 2693 27 2707
rect 53 2693 67 2707
rect 53 2653 67 2667
rect 33 2573 47 2587
rect 13 2553 27 2567
rect 173 2933 187 2947
rect 233 3113 247 3127
rect 413 3673 427 3687
rect 373 3653 387 3667
rect 493 3713 507 3727
rect 513 3733 527 3747
rect 593 3753 607 3767
rect 633 3753 647 3767
rect 573 3713 587 3727
rect 513 3693 527 3707
rect 533 3693 547 3707
rect 573 3693 587 3707
rect 513 3653 527 3667
rect 433 3633 447 3647
rect 453 3633 467 3647
rect 373 3613 387 3627
rect 333 3573 347 3587
rect 353 3573 367 3587
rect 533 3573 547 3587
rect 373 3493 387 3507
rect 373 3453 387 3467
rect 513 3533 527 3547
rect 473 3513 487 3527
rect 433 3493 447 3507
rect 493 3493 507 3507
rect 533 3493 547 3507
rect 553 3513 567 3527
rect 553 3473 567 3487
rect 413 3453 427 3467
rect 313 3313 327 3327
rect 293 3273 307 3287
rect 333 3273 347 3287
rect 533 3353 547 3367
rect 393 3313 407 3327
rect 453 3313 467 3327
rect 453 3293 467 3307
rect 513 3313 527 3327
rect 393 3273 407 3287
rect 373 3233 387 3247
rect 413 3233 427 3247
rect 433 3253 447 3267
rect 353 3213 367 3227
rect 433 3213 447 3227
rect 353 3193 367 3207
rect 313 3173 327 3187
rect 333 3173 347 3187
rect 293 3133 307 3147
rect 273 3113 287 3127
rect 253 3073 267 3087
rect 213 2993 227 3007
rect 193 2853 207 2867
rect 133 2773 147 2787
rect 153 2773 167 2787
rect 293 3013 307 3027
rect 293 2993 307 3007
rect 253 2893 267 2907
rect 233 2813 247 2827
rect 273 2813 287 2827
rect 213 2773 227 2787
rect 113 2733 127 2747
rect 173 2733 187 2747
rect 193 2753 207 2767
rect 233 2753 247 2767
rect 373 3173 387 3187
rect 393 3153 407 3167
rect 313 2913 327 2927
rect 373 3033 387 3047
rect 373 2993 387 3007
rect 373 2953 387 2967
rect 473 3253 487 3267
rect 473 3213 487 3227
rect 453 3173 467 3187
rect 453 3153 467 3167
rect 433 3113 447 3127
rect 433 2953 447 2967
rect 353 2873 367 2887
rect 333 2793 347 2807
rect 293 2773 307 2787
rect 353 2773 367 2787
rect 373 2773 387 2787
rect 253 2733 267 2747
rect 273 2733 287 2747
rect 93 2653 107 2667
rect 93 2613 107 2627
rect 73 2553 87 2567
rect 53 2533 67 2547
rect 13 2493 27 2507
rect 33 2393 47 2407
rect 193 2713 207 2727
rect 293 2713 307 2727
rect 213 2693 227 2707
rect 173 2613 187 2627
rect 153 2593 167 2607
rect 133 2573 147 2587
rect 113 2533 127 2547
rect 153 2533 167 2547
rect 13 2313 27 2327
rect 33 2313 47 2327
rect 93 2313 107 2327
rect 53 2273 67 2287
rect 93 2273 107 2287
rect 33 2253 47 2267
rect 13 2173 27 2187
rect 73 2253 87 2267
rect 53 2093 67 2107
rect 73 2093 87 2107
rect 53 2073 67 2087
rect 13 1993 27 2007
rect 13 1873 27 1887
rect 33 1853 47 1867
rect 133 2353 147 2367
rect 253 2593 267 2607
rect 393 2753 407 2767
rect 373 2733 387 2747
rect 353 2713 367 2727
rect 413 2733 427 2747
rect 433 2733 447 2747
rect 333 2693 347 2707
rect 313 2653 327 2667
rect 233 2533 247 2547
rect 253 2533 267 2547
rect 213 2393 227 2407
rect 193 2293 207 2307
rect 313 2513 327 2527
rect 353 2613 367 2627
rect 413 2653 427 2667
rect 433 2613 447 2627
rect 473 3093 487 3107
rect 513 3073 527 3087
rect 553 3293 567 3307
rect 553 3193 567 3207
rect 813 4173 827 4187
rect 853 4173 867 4187
rect 913 4413 927 4427
rect 1053 4393 1067 4407
rect 1093 4453 1107 4467
rect 1153 4473 1167 4487
rect 1173 4473 1187 4487
rect 1133 4433 1147 4447
rect 1293 4533 1307 4547
rect 1453 4533 1467 4547
rect 1273 4493 1287 4507
rect 1433 4513 1447 4527
rect 1313 4493 1327 4507
rect 1353 4493 1367 4507
rect 1193 4453 1207 4467
rect 1093 4413 1107 4427
rect 1173 4413 1187 4427
rect 913 4353 927 4367
rect 953 4353 967 4367
rect 1073 4353 1087 4367
rect 1153 4353 1167 4367
rect 913 4213 927 4227
rect 893 4173 907 4187
rect 953 4193 967 4207
rect 1053 4213 1067 4227
rect 873 4153 887 4167
rect 933 4153 947 4167
rect 773 4133 787 4147
rect 893 4133 907 4147
rect 1033 4133 1047 4147
rect 713 4013 727 4027
rect 793 4053 807 4067
rect 773 3993 787 4007
rect 853 4033 867 4047
rect 753 3973 767 3987
rect 773 3953 787 3967
rect 813 3973 827 3987
rect 753 3933 767 3947
rect 833 3953 847 3967
rect 933 4033 947 4047
rect 953 4033 967 4047
rect 1113 4213 1127 4227
rect 1093 4173 1107 4187
rect 1073 4113 1087 4127
rect 1073 4053 1087 4067
rect 973 3973 987 3987
rect 993 3993 1007 4007
rect 1013 3993 1027 4007
rect 1033 3973 1047 3987
rect 973 3953 987 3967
rect 873 3933 887 3947
rect 693 3913 707 3927
rect 853 3913 867 3927
rect 833 3773 847 3787
rect 673 3693 687 3707
rect 693 3713 707 3727
rect 733 3713 747 3727
rect 793 3713 807 3727
rect 753 3693 767 3707
rect 593 3573 607 3587
rect 653 3593 667 3607
rect 693 3673 707 3687
rect 833 3673 847 3687
rect 793 3633 807 3647
rect 693 3613 707 3627
rect 753 3613 767 3627
rect 673 3553 687 3567
rect 733 3553 747 3567
rect 653 3513 667 3527
rect 613 3393 627 3407
rect 593 3293 607 3307
rect 593 3253 607 3267
rect 593 3213 607 3227
rect 593 3173 607 3187
rect 573 3153 587 3167
rect 693 3493 707 3507
rect 673 3453 687 3467
rect 693 3453 707 3467
rect 673 3353 687 3367
rect 633 3333 647 3347
rect 653 3253 667 3267
rect 653 3173 667 3187
rect 613 3153 627 3167
rect 653 3153 667 3167
rect 633 3133 647 3147
rect 553 3093 567 3107
rect 573 3093 587 3107
rect 593 3093 607 3107
rect 533 3053 547 3067
rect 513 3033 527 3047
rect 533 3013 547 3027
rect 473 2973 487 2987
rect 453 2573 467 2587
rect 393 2553 407 2567
rect 413 2533 427 2547
rect 433 2533 447 2547
rect 353 2513 367 2527
rect 373 2513 387 2527
rect 333 2453 347 2467
rect 273 2353 287 2367
rect 313 2353 327 2367
rect 413 2413 427 2427
rect 413 2333 427 2347
rect 313 2313 327 2327
rect 353 2313 367 2327
rect 293 2293 307 2307
rect 133 2253 147 2267
rect 173 2273 187 2287
rect 233 2273 247 2287
rect 273 2273 287 2287
rect 193 2233 207 2247
rect 213 2233 227 2247
rect 213 2213 227 2227
rect 233 2213 247 2227
rect 153 2193 167 2207
rect 173 2133 187 2147
rect 313 2273 327 2287
rect 353 2273 367 2287
rect 333 2253 347 2267
rect 373 2253 387 2267
rect 293 2233 307 2247
rect 333 2233 347 2247
rect 273 2213 287 2227
rect 353 2193 367 2207
rect 313 2173 327 2187
rect 273 2153 287 2167
rect 133 2073 147 2087
rect 173 2073 187 2087
rect 213 2073 227 2087
rect 233 2073 247 2087
rect 253 2073 267 2087
rect 353 2093 367 2107
rect 73 2033 87 2047
rect 93 2033 107 2047
rect 53 1833 67 1847
rect 93 1873 107 1887
rect 113 1833 127 1847
rect 73 1813 87 1827
rect 93 1813 107 1827
rect 173 2033 187 2047
rect 273 2053 287 2067
rect 293 2053 307 2067
rect 313 2053 327 2067
rect 353 2073 367 2087
rect 253 2033 267 2047
rect 173 1973 187 1987
rect 233 2013 247 2027
rect 213 1953 227 1967
rect 233 1933 247 1947
rect 293 1933 307 1947
rect 233 1913 247 1927
rect 213 1853 227 1867
rect 333 2033 347 2047
rect 313 1893 327 1907
rect 293 1853 307 1867
rect 233 1833 247 1847
rect 213 1813 227 1827
rect 73 1773 87 1787
rect 153 1793 167 1807
rect 193 1793 207 1807
rect 93 1753 107 1767
rect 33 1733 47 1747
rect 13 1713 27 1727
rect 173 1733 187 1747
rect 133 1713 147 1727
rect 113 1693 127 1707
rect 133 1673 147 1687
rect 13 1593 27 1607
rect 33 1573 47 1587
rect 93 1613 107 1627
rect 133 1613 147 1627
rect 173 1613 187 1627
rect 93 1593 107 1607
rect 113 1573 127 1587
rect 133 1573 147 1587
rect 153 1573 167 1587
rect 113 1553 127 1567
rect 53 1393 67 1407
rect 73 1393 87 1407
rect 253 1793 267 1807
rect 273 1773 287 1787
rect 253 1753 267 1767
rect 213 1733 227 1747
rect 253 1693 267 1707
rect 273 1693 287 1707
rect 213 1573 227 1587
rect 193 1553 207 1567
rect 273 1633 287 1647
rect 453 2513 467 2527
rect 493 2933 507 2947
rect 593 3073 607 3087
rect 593 3033 607 3047
rect 573 2993 587 3007
rect 593 3013 607 3027
rect 613 2933 627 2947
rect 553 2913 567 2927
rect 573 2893 587 2907
rect 553 2833 567 2847
rect 553 2813 567 2827
rect 533 2793 547 2807
rect 713 3373 727 3387
rect 753 3533 767 3547
rect 833 3533 847 3547
rect 833 3513 847 3527
rect 753 3373 767 3387
rect 733 3353 747 3367
rect 813 3433 827 3447
rect 773 3333 787 3347
rect 793 3273 807 3287
rect 733 3213 747 3227
rect 733 3193 747 3207
rect 873 3793 887 3807
rect 953 3773 967 3787
rect 913 3733 927 3747
rect 1093 3953 1107 3967
rect 1033 3933 1047 3947
rect 1273 4453 1287 4467
rect 1333 4473 1347 4487
rect 1253 4433 1267 4447
rect 1453 4493 1467 4507
rect 1393 4473 1407 4487
rect 1373 4453 1387 4467
rect 1353 4413 1367 4427
rect 1633 4533 1647 4547
rect 2273 4533 2287 4547
rect 2333 4533 2347 4547
rect 3333 4533 3347 4547
rect 3433 4533 3447 4547
rect 3953 4533 3967 4547
rect 1613 4513 1627 4527
rect 1553 4493 1567 4507
rect 1493 4473 1507 4487
rect 1573 4473 1587 4487
rect 1553 4453 1567 4467
rect 1593 4453 1607 4467
rect 1513 4433 1527 4447
rect 1693 4513 1707 4527
rect 1813 4513 1827 4527
rect 1953 4513 1967 4527
rect 2013 4513 2027 4527
rect 2053 4513 2067 4527
rect 1653 4453 1667 4467
rect 1773 4493 1787 4507
rect 1693 4433 1707 4447
rect 1593 4413 1607 4427
rect 1253 4393 1267 4407
rect 1413 4393 1427 4407
rect 1553 4393 1567 4407
rect 1213 4373 1227 4387
rect 1673 4253 1687 4267
rect 1393 4233 1407 4247
rect 1553 4233 1567 4247
rect 1233 4193 1247 4207
rect 1293 4213 1307 4227
rect 1313 4193 1327 4207
rect 1433 4213 1447 4227
rect 1473 4213 1487 4227
rect 1453 4193 1467 4207
rect 1233 4173 1247 4187
rect 1273 4173 1287 4187
rect 1333 4173 1347 4187
rect 1133 4133 1147 4147
rect 1193 4133 1207 4147
rect 1213 4033 1227 4047
rect 1133 3973 1147 3987
rect 1113 3893 1127 3907
rect 1333 4113 1347 4127
rect 1233 4013 1247 4027
rect 1193 3953 1207 3967
rect 1393 4173 1407 4187
rect 1353 4093 1367 4107
rect 1373 4033 1387 4047
rect 1353 4013 1367 4027
rect 1293 3973 1307 3987
rect 1333 3973 1347 3987
rect 1453 4133 1467 4147
rect 1413 4113 1427 4127
rect 1413 4093 1427 4107
rect 1393 3993 1407 4007
rect 1393 3953 1407 3967
rect 1433 4013 1447 4027
rect 1493 4153 1507 4167
rect 1913 4493 1927 4507
rect 1893 4453 1907 4467
rect 1993 4473 2007 4487
rect 2013 4453 2027 4467
rect 2173 4493 2187 4507
rect 1753 4393 1767 4407
rect 1833 4433 1847 4447
rect 1973 4433 1987 4447
rect 2033 4393 2047 4407
rect 1793 4313 1807 4327
rect 1893 4313 1907 4327
rect 1933 4313 1947 4327
rect 1793 4233 1807 4247
rect 1553 4193 1567 4207
rect 1533 4073 1547 4087
rect 1473 4013 1487 4027
rect 1513 3993 1527 4007
rect 1453 3953 1467 3967
rect 1493 3953 1507 3967
rect 1413 3933 1427 3947
rect 1473 3933 1487 3947
rect 1233 3893 1247 3907
rect 1273 3893 1287 3907
rect 1033 3793 1047 3807
rect 1173 3793 1187 3807
rect 993 3753 1007 3767
rect 1033 3733 1047 3747
rect 1073 3733 1087 3747
rect 973 3713 987 3727
rect 933 3693 947 3707
rect 1053 3713 1067 3727
rect 1013 3693 1027 3707
rect 1053 3693 1067 3707
rect 1093 3713 1107 3727
rect 1113 3733 1127 3747
rect 913 3673 927 3687
rect 933 3673 947 3687
rect 973 3673 987 3687
rect 1073 3673 1087 3687
rect 873 3533 887 3547
rect 873 3493 887 3507
rect 893 3493 907 3507
rect 853 3393 867 3407
rect 833 3293 847 3307
rect 813 3253 827 3267
rect 933 3653 947 3667
rect 1073 3633 1087 3647
rect 1133 3693 1147 3707
rect 1193 3713 1207 3727
rect 1173 3673 1187 3687
rect 1213 3673 1227 3687
rect 1133 3613 1147 3627
rect 1073 3593 1087 3607
rect 1093 3593 1107 3607
rect 993 3573 1007 3587
rect 1113 3573 1127 3587
rect 973 3553 987 3567
rect 1013 3533 1027 3547
rect 1053 3533 1067 3547
rect 1093 3533 1107 3547
rect 993 3513 1007 3527
rect 1013 3493 1027 3507
rect 1033 3493 1047 3507
rect 1153 3573 1167 3587
rect 1333 3853 1347 3867
rect 1413 3753 1427 3767
rect 1273 3713 1287 3727
rect 1373 3733 1387 3747
rect 1353 3713 1367 3727
rect 1433 3713 1447 3727
rect 1733 4193 1747 4207
rect 1833 4213 1847 4227
rect 1813 4193 1827 4207
rect 1873 4213 1887 4227
rect 1933 4233 1947 4247
rect 1913 4213 1927 4227
rect 1893 4193 1907 4207
rect 1973 4213 1987 4227
rect 2013 4213 2027 4227
rect 1753 4173 1767 4187
rect 1673 4153 1687 4167
rect 1613 4093 1627 4107
rect 1653 4093 1667 4107
rect 1653 4013 1667 4027
rect 1593 3993 1607 4007
rect 1633 3993 1647 4007
rect 1713 4113 1727 4127
rect 1713 4093 1727 4107
rect 1933 4173 1947 4187
rect 1893 4153 1907 4167
rect 1853 4133 1867 4147
rect 1873 4073 1887 4087
rect 1813 4053 1827 4067
rect 1793 4033 1807 4047
rect 1673 3993 1687 4007
rect 1693 3993 1707 4007
rect 1753 3993 1767 4007
rect 1773 3993 1787 4007
rect 1533 3933 1547 3947
rect 1513 3853 1527 3867
rect 1573 3853 1587 3867
rect 1633 3753 1647 3767
rect 1573 3733 1587 3747
rect 1493 3713 1507 3727
rect 1473 3693 1487 3707
rect 1513 3693 1527 3707
rect 1533 3713 1547 3727
rect 1553 3693 1567 3707
rect 1253 3673 1267 3687
rect 1393 3673 1407 3687
rect 1413 3673 1427 3687
rect 1453 3673 1467 3687
rect 1253 3653 1267 3667
rect 1373 3633 1387 3647
rect 1273 3553 1287 3567
rect 1233 3533 1247 3547
rect 1113 3493 1127 3507
rect 1153 3493 1167 3507
rect 993 3473 1007 3487
rect 1033 3473 1047 3487
rect 1093 3473 1107 3487
rect 1073 3433 1087 3447
rect 933 3393 947 3407
rect 1013 3393 1027 3407
rect 913 3353 927 3367
rect 973 3353 987 3367
rect 913 3273 927 3287
rect 873 3253 887 3267
rect 853 3213 867 3227
rect 873 3233 887 3247
rect 933 3233 947 3247
rect 953 3253 967 3267
rect 893 3213 907 3227
rect 673 3133 687 3147
rect 673 2993 687 3007
rect 693 3013 707 3027
rect 713 2993 727 3007
rect 673 2973 687 2987
rect 653 2893 667 2907
rect 613 2833 627 2847
rect 573 2773 587 2787
rect 493 2753 507 2767
rect 493 2733 507 2747
rect 553 2733 567 2747
rect 573 2733 587 2747
rect 533 2713 547 2727
rect 513 2573 527 2587
rect 553 2593 567 2607
rect 533 2533 547 2547
rect 533 2513 547 2527
rect 473 2473 487 2487
rect 613 2733 627 2747
rect 693 2953 707 2967
rect 713 2953 727 2967
rect 673 2813 687 2827
rect 793 3193 807 3207
rect 813 3193 827 3207
rect 833 3193 847 3207
rect 773 3173 787 3187
rect 753 3153 767 3167
rect 793 3093 807 3107
rect 753 3033 767 3047
rect 873 3173 887 3187
rect 873 3153 887 3167
rect 833 3053 847 3067
rect 833 3033 847 3047
rect 853 3033 867 3047
rect 813 2993 827 3007
rect 773 2973 787 2987
rect 753 2933 767 2947
rect 733 2833 747 2847
rect 713 2793 727 2807
rect 753 2793 767 2807
rect 993 3273 1007 3287
rect 1093 3373 1107 3387
rect 1093 3333 1107 3347
rect 1133 3333 1147 3347
rect 993 3233 1007 3247
rect 1053 3253 1067 3267
rect 1073 3233 1087 3247
rect 1073 3213 1087 3227
rect 933 3153 947 3167
rect 973 3153 987 3167
rect 913 3113 927 3127
rect 993 3093 1007 3107
rect 1073 3093 1087 3107
rect 973 3033 987 3047
rect 933 2993 947 3007
rect 893 2973 907 2987
rect 873 2953 887 2967
rect 873 2893 887 2907
rect 853 2833 867 2847
rect 833 2813 847 2827
rect 673 2733 687 2747
rect 613 2693 627 2707
rect 653 2693 667 2707
rect 613 2613 627 2627
rect 593 2593 607 2607
rect 613 2573 627 2587
rect 733 2733 747 2747
rect 813 2773 827 2787
rect 833 2753 847 2767
rect 773 2693 787 2707
rect 713 2573 727 2587
rect 613 2513 627 2527
rect 573 2493 587 2507
rect 593 2473 607 2487
rect 493 2413 507 2427
rect 573 2413 587 2427
rect 453 2353 467 2367
rect 513 2313 527 2327
rect 433 2273 447 2287
rect 473 2253 487 2267
rect 433 2233 447 2247
rect 473 2233 487 2247
rect 393 2213 407 2227
rect 453 2113 467 2127
rect 473 2093 487 2107
rect 393 2053 407 2067
rect 413 2053 427 2067
rect 433 2053 447 2067
rect 533 2273 547 2287
rect 553 2253 567 2267
rect 513 2213 527 2227
rect 393 2033 407 2047
rect 393 1873 407 1887
rect 373 1853 387 1867
rect 433 2033 447 2047
rect 453 1853 467 1867
rect 413 1833 427 1847
rect 333 1813 347 1827
rect 373 1813 387 1827
rect 433 1813 447 1827
rect 593 2253 607 2267
rect 813 2733 827 2747
rect 853 2733 867 2747
rect 813 2653 827 2667
rect 833 2653 847 2667
rect 793 2633 807 2647
rect 793 2613 807 2627
rect 693 2513 707 2527
rect 673 2373 687 2387
rect 753 2513 767 2527
rect 713 2473 727 2487
rect 853 2613 867 2627
rect 833 2553 847 2567
rect 893 2833 907 2847
rect 893 2733 907 2747
rect 913 2733 927 2747
rect 1033 3073 1047 3087
rect 1013 3053 1027 3067
rect 1133 3293 1147 3307
rect 1113 3213 1127 3227
rect 1133 3153 1147 3167
rect 1113 3133 1127 3147
rect 1193 3473 1207 3487
rect 1233 3493 1247 3507
rect 1253 3473 1267 3487
rect 1253 3413 1267 3427
rect 1213 3393 1227 3407
rect 1213 3313 1227 3327
rect 1173 3293 1187 3307
rect 1293 3473 1307 3487
rect 1313 3493 1327 3507
rect 1413 3513 1427 3527
rect 1433 3493 1447 3507
rect 1333 3473 1347 3487
rect 1373 3473 1387 3487
rect 1373 3353 1387 3367
rect 1173 3253 1187 3267
rect 1173 3193 1187 3207
rect 1173 3093 1187 3107
rect 1253 3253 1267 3267
rect 1273 3253 1287 3267
rect 1273 3233 1287 3247
rect 1213 3153 1227 3167
rect 1233 3153 1247 3167
rect 1213 3113 1227 3127
rect 1193 3073 1207 3087
rect 1153 3053 1167 3067
rect 1173 3053 1187 3067
rect 993 2993 1007 3007
rect 1013 2953 1027 2967
rect 1053 2953 1067 2967
rect 953 2933 967 2947
rect 953 2773 967 2787
rect 933 2633 947 2647
rect 913 2573 927 2587
rect 893 2553 907 2567
rect 833 2513 847 2527
rect 873 2533 887 2547
rect 1253 3073 1267 3087
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1333 3193 1347 3207
rect 1433 3333 1447 3347
rect 1393 3253 1407 3267
rect 1433 3213 1447 3227
rect 1413 3153 1427 3167
rect 1393 3133 1407 3147
rect 1293 3073 1307 3087
rect 1173 3013 1187 3027
rect 1233 3013 1247 3027
rect 1273 3033 1287 3047
rect 1093 2933 1107 2947
rect 1253 2993 1267 3007
rect 1273 2993 1287 3007
rect 1593 3713 1607 3727
rect 1673 3713 1687 3727
rect 1573 3673 1587 3687
rect 1613 3673 1627 3687
rect 1753 3713 1767 3727
rect 1693 3693 1707 3707
rect 1713 3693 1727 3707
rect 1733 3693 1747 3707
rect 1653 3673 1667 3687
rect 1773 3693 1787 3707
rect 1753 3673 1767 3687
rect 1553 3653 1567 3667
rect 1633 3633 1647 3647
rect 1573 3613 1587 3627
rect 1533 3593 1547 3607
rect 1553 3513 1567 3527
rect 1473 3393 1487 3407
rect 1453 3193 1467 3207
rect 1493 3253 1507 3267
rect 1513 3253 1527 3267
rect 1553 3233 1567 3247
rect 1533 3213 1547 3227
rect 1553 3193 1567 3207
rect 1493 3173 1507 3187
rect 1513 3173 1527 3187
rect 1473 3153 1487 3167
rect 1493 3093 1507 3107
rect 1473 3073 1487 3087
rect 1513 3073 1527 3087
rect 1233 2973 1247 2987
rect 1113 2873 1127 2887
rect 1173 2873 1187 2887
rect 1053 2813 1067 2827
rect 973 2733 987 2747
rect 1013 2753 1027 2767
rect 1093 2773 1107 2787
rect 1053 2733 1067 2747
rect 1073 2733 1087 2747
rect 973 2653 987 2667
rect 953 2593 967 2607
rect 1013 2713 1027 2727
rect 993 2633 1007 2647
rect 953 2573 967 2587
rect 973 2573 987 2587
rect 1033 2693 1047 2707
rect 1033 2613 1047 2627
rect 873 2513 887 2527
rect 993 2553 1007 2567
rect 1013 2553 1027 2567
rect 1133 2813 1147 2827
rect 1113 2693 1127 2707
rect 1193 2793 1207 2807
rect 1193 2773 1207 2787
rect 1153 2733 1167 2747
rect 1173 2733 1187 2747
rect 1293 2953 1307 2967
rect 1253 2773 1267 2787
rect 1213 2693 1227 2707
rect 1133 2673 1147 2687
rect 1093 2653 1107 2667
rect 1253 2693 1267 2707
rect 1353 2873 1367 2887
rect 1313 2813 1327 2827
rect 1293 2713 1307 2727
rect 1133 2633 1147 2647
rect 1153 2633 1167 2647
rect 1233 2633 1247 2647
rect 1093 2593 1107 2607
rect 1053 2553 1067 2567
rect 953 2513 967 2527
rect 933 2493 947 2507
rect 813 2473 827 2487
rect 833 2473 847 2487
rect 773 2453 787 2467
rect 753 2393 767 2407
rect 633 2313 647 2327
rect 653 2293 667 2307
rect 753 2353 767 2367
rect 733 2293 747 2307
rect 673 2273 687 2287
rect 693 2273 707 2287
rect 573 2213 587 2227
rect 553 2193 567 2207
rect 533 2153 547 2167
rect 673 2213 687 2227
rect 653 2193 667 2207
rect 573 2173 587 2187
rect 573 2113 587 2127
rect 513 2033 527 2047
rect 553 2033 567 2047
rect 513 1993 527 2007
rect 473 1833 487 1847
rect 333 1773 347 1787
rect 313 1713 327 1727
rect 293 1613 307 1627
rect 293 1573 307 1587
rect 193 1453 207 1467
rect 93 1373 107 1387
rect 133 1373 147 1387
rect 53 1333 67 1347
rect 233 1373 247 1387
rect 313 1533 327 1547
rect 293 1433 307 1447
rect 253 1353 267 1367
rect 273 1353 287 1367
rect 373 1773 387 1787
rect 453 1773 467 1787
rect 493 1773 507 1787
rect 353 1753 367 1767
rect 353 1653 367 1667
rect 553 1913 567 1927
rect 533 1773 547 1787
rect 593 2053 607 2067
rect 633 2113 647 2127
rect 653 2073 667 2087
rect 633 2053 647 2067
rect 633 2013 647 2027
rect 613 1893 627 1907
rect 573 1853 587 1867
rect 573 1813 587 1827
rect 613 1773 627 1787
rect 653 1973 667 1987
rect 713 2173 727 2187
rect 753 2133 767 2147
rect 713 2113 727 2127
rect 813 2393 827 2407
rect 793 2253 807 2267
rect 913 2453 927 2467
rect 873 2393 887 2407
rect 913 2293 927 2307
rect 853 2253 867 2267
rect 833 2233 847 2247
rect 833 2213 847 2227
rect 813 2193 827 2207
rect 793 2113 807 2127
rect 773 2093 787 2107
rect 793 2093 807 2107
rect 693 2053 707 2067
rect 713 2033 727 2047
rect 693 1953 707 1967
rect 673 1913 687 1927
rect 753 2033 767 2047
rect 733 1993 747 2007
rect 713 1893 727 1907
rect 713 1833 727 1847
rect 673 1813 687 1827
rect 673 1793 687 1807
rect 693 1773 707 1787
rect 533 1753 547 1767
rect 593 1753 607 1767
rect 633 1753 647 1767
rect 413 1733 427 1747
rect 513 1733 527 1747
rect 393 1713 407 1727
rect 453 1693 467 1707
rect 413 1633 427 1647
rect 373 1593 387 1607
rect 373 1573 387 1587
rect 413 1573 427 1587
rect 433 1593 447 1607
rect 433 1553 447 1567
rect 373 1433 387 1447
rect 353 1413 367 1427
rect 353 1393 367 1407
rect 93 1313 107 1327
rect 113 1313 127 1327
rect 13 1133 27 1147
rect 173 1333 187 1347
rect 233 1333 247 1347
rect 153 1293 167 1307
rect 173 1293 187 1307
rect 73 1273 87 1287
rect 133 1273 147 1287
rect 53 1253 67 1267
rect 153 1153 167 1167
rect 93 1133 107 1147
rect 113 1133 127 1147
rect 13 1113 27 1127
rect 33 1113 47 1127
rect 33 1093 47 1107
rect 73 1093 87 1107
rect 133 1093 147 1107
rect 173 1113 187 1127
rect 213 1173 227 1187
rect 253 1313 267 1327
rect 233 1133 247 1147
rect 213 1113 227 1127
rect 93 1073 107 1087
rect 13 933 27 947
rect 73 873 87 887
rect 13 793 27 807
rect 353 1353 367 1367
rect 413 1413 427 1427
rect 393 1373 407 1387
rect 493 1633 507 1647
rect 473 1613 487 1627
rect 473 1493 487 1507
rect 453 1453 467 1467
rect 433 1393 447 1407
rect 333 1333 347 1347
rect 353 1313 367 1327
rect 393 1333 407 1347
rect 413 1333 427 1347
rect 653 1733 667 1747
rect 653 1713 667 1727
rect 633 1653 647 1667
rect 573 1633 587 1647
rect 593 1633 607 1647
rect 533 1613 547 1627
rect 633 1613 647 1627
rect 733 1813 747 1827
rect 733 1773 747 1787
rect 913 2253 927 2267
rect 993 2513 1007 2527
rect 1073 2513 1087 2527
rect 973 2493 987 2507
rect 953 2473 967 2487
rect 973 2433 987 2447
rect 953 2333 967 2347
rect 953 2293 967 2307
rect 953 2253 967 2267
rect 1013 2473 1027 2487
rect 1033 2393 1047 2407
rect 993 2373 1007 2387
rect 993 2293 1007 2307
rect 1033 2273 1047 2287
rect 1073 2433 1087 2447
rect 1173 2593 1187 2607
rect 1233 2593 1247 2607
rect 1193 2573 1207 2587
rect 1233 2573 1247 2587
rect 1153 2533 1167 2547
rect 1153 2513 1167 2527
rect 1193 2513 1207 2527
rect 1133 2493 1147 2507
rect 1113 2453 1127 2467
rect 1153 2373 1167 2387
rect 1113 2313 1127 2327
rect 1133 2313 1147 2327
rect 1093 2293 1107 2307
rect 1013 2253 1027 2267
rect 1053 2253 1067 2267
rect 1073 2253 1087 2267
rect 1413 2993 1427 3007
rect 1593 3553 1607 3567
rect 1593 3473 1607 3487
rect 1813 4013 1827 4027
rect 1973 4153 1987 4167
rect 1933 4033 1947 4047
rect 1913 4013 1927 4027
rect 1833 3993 1847 4007
rect 1953 4013 1967 4027
rect 1913 3973 1927 3987
rect 1833 3953 1847 3967
rect 1853 3953 1867 3967
rect 1813 3933 1827 3947
rect 1893 3753 1907 3767
rect 1813 3693 1827 3707
rect 1993 4093 2007 4107
rect 2133 4453 2147 4467
rect 2193 4453 2207 4467
rect 2213 4473 2227 4487
rect 2253 4433 2267 4447
rect 2093 4313 2107 4327
rect 2113 4273 2127 4287
rect 2093 4193 2107 4207
rect 2073 4133 2087 4147
rect 2293 4513 2307 4527
rect 2393 4493 2407 4507
rect 2473 4493 2487 4507
rect 2513 4493 2527 4507
rect 2313 4453 2327 4467
rect 2373 4473 2387 4487
rect 2433 4473 2447 4487
rect 2353 4433 2367 4447
rect 2133 4113 2147 4127
rect 2173 4113 2187 4127
rect 2073 4093 2087 4107
rect 2053 4033 2067 4047
rect 1973 3973 1987 3987
rect 2093 3973 2107 3987
rect 2153 3973 2167 3987
rect 1993 3953 2007 3967
rect 2353 4173 2367 4187
rect 2313 4093 2327 4107
rect 2273 4073 2287 4087
rect 2253 4053 2267 4067
rect 2213 3973 2227 3987
rect 2273 4033 2287 4047
rect 2273 3993 2287 4007
rect 2453 4453 2467 4467
rect 2493 4433 2507 4447
rect 2533 4433 2547 4447
rect 2433 4413 2447 4427
rect 2413 4393 2427 4407
rect 2373 4033 2387 4047
rect 2393 4013 2407 4027
rect 2453 4373 2467 4387
rect 2613 4473 2627 4487
rect 2653 4473 2667 4487
rect 2713 4453 2727 4467
rect 2673 4433 2687 4447
rect 2573 4413 2587 4427
rect 2633 4413 2647 4427
rect 2793 4473 2807 4487
rect 2673 4233 2687 4247
rect 2493 4193 2507 4207
rect 2553 4173 2567 4187
rect 2593 4173 2607 4187
rect 2633 4173 2647 4187
rect 2513 4153 2527 4167
rect 2553 4153 2567 4167
rect 2593 4153 2607 4167
rect 2433 4013 2447 4027
rect 2573 4013 2587 4027
rect 2353 3993 2367 4007
rect 1953 3753 1967 3767
rect 1933 3733 1947 3747
rect 1973 3733 1987 3747
rect 1953 3693 1967 3707
rect 2053 3713 2067 3727
rect 1873 3673 1887 3687
rect 1913 3673 1927 3687
rect 1953 3673 1967 3687
rect 1993 3673 2007 3687
rect 1833 3653 1847 3667
rect 1693 3533 1707 3547
rect 1793 3533 1807 3547
rect 1833 3533 1847 3547
rect 1673 3513 1687 3527
rect 1673 3473 1687 3487
rect 1673 3413 1687 3427
rect 1673 3373 1687 3387
rect 1633 3313 1647 3327
rect 1593 3253 1607 3267
rect 1613 3233 1627 3247
rect 1633 3253 1647 3267
rect 1713 3513 1727 3527
rect 1793 3513 1807 3527
rect 1753 3493 1767 3507
rect 1853 3493 1867 3507
rect 1733 3453 1747 3467
rect 1753 3453 1767 3467
rect 1713 3393 1727 3407
rect 1713 3353 1727 3367
rect 1733 3353 1747 3367
rect 1693 3253 1707 3267
rect 1613 3153 1627 3167
rect 1573 3033 1587 3047
rect 1473 2993 1487 3007
rect 1513 3013 1527 3027
rect 1553 3013 1567 3027
rect 1553 2993 1567 3007
rect 1393 2973 1407 2987
rect 1373 2793 1387 2807
rect 1353 2753 1367 2767
rect 1313 2653 1327 2667
rect 1333 2653 1347 2667
rect 1293 2613 1307 2627
rect 1333 2593 1347 2607
rect 1373 2733 1387 2747
rect 1373 2573 1387 2587
rect 1273 2553 1287 2567
rect 1353 2553 1367 2567
rect 1273 2493 1287 2507
rect 1253 2393 1267 2407
rect 1193 2333 1207 2347
rect 1253 2293 1267 2307
rect 1173 2273 1187 2287
rect 1173 2253 1187 2267
rect 1213 2273 1227 2287
rect 1233 2253 1247 2267
rect 953 2233 967 2247
rect 973 2233 987 2247
rect 1093 2233 1107 2247
rect 933 2213 947 2227
rect 913 2193 927 2207
rect 893 2153 907 2167
rect 933 2113 947 2127
rect 893 2093 907 2107
rect 813 2073 827 2087
rect 973 2213 987 2227
rect 1133 2213 1147 2227
rect 1153 2213 1167 2227
rect 813 2053 827 2067
rect 933 2073 947 2087
rect 953 2073 967 2087
rect 913 2053 927 2067
rect 793 2013 807 2027
rect 873 2033 887 2047
rect 913 2033 927 2047
rect 773 1993 787 2007
rect 853 1993 867 2007
rect 853 1953 867 1967
rect 773 1913 787 1927
rect 833 1873 847 1887
rect 813 1853 827 1867
rect 813 1813 827 1827
rect 893 2013 907 2027
rect 933 2013 947 2027
rect 893 1973 907 1987
rect 893 1873 907 1887
rect 873 1853 887 1867
rect 853 1833 867 1847
rect 1033 2113 1047 2127
rect 1013 2093 1027 2107
rect 993 2073 1007 2087
rect 1113 2093 1127 2107
rect 1153 2073 1167 2087
rect 1013 2053 1027 2067
rect 1013 2033 1027 2047
rect 1093 2053 1107 2067
rect 1133 2053 1147 2067
rect 1153 2033 1167 2047
rect 993 2013 1007 2027
rect 1033 2013 1047 2027
rect 1053 2013 1067 2027
rect 1093 2013 1107 2027
rect 973 1993 987 2007
rect 993 1973 1007 1987
rect 1013 1893 1027 1907
rect 953 1873 967 1887
rect 953 1853 967 1867
rect 913 1813 927 1827
rect 793 1793 807 1807
rect 753 1733 767 1747
rect 753 1693 767 1707
rect 713 1633 727 1647
rect 653 1593 667 1607
rect 573 1573 587 1587
rect 613 1573 627 1587
rect 333 1293 347 1307
rect 373 1293 387 1307
rect 413 1313 427 1327
rect 533 1533 547 1547
rect 553 1513 567 1527
rect 493 1313 507 1327
rect 513 1313 527 1327
rect 533 1313 547 1327
rect 313 1273 327 1287
rect 273 1213 287 1227
rect 293 1193 307 1207
rect 353 1273 367 1287
rect 293 1173 307 1187
rect 333 1173 347 1187
rect 373 1173 387 1187
rect 433 1233 447 1247
rect 453 1213 467 1227
rect 493 1273 507 1287
rect 553 1273 567 1287
rect 373 1153 387 1167
rect 393 1153 407 1167
rect 413 1153 427 1167
rect 333 1133 347 1147
rect 353 1133 367 1147
rect 253 1113 267 1127
rect 293 1113 307 1127
rect 253 1093 267 1107
rect 373 1113 387 1127
rect 273 1073 287 1087
rect 173 1053 187 1067
rect 193 1053 207 1067
rect 253 1053 267 1067
rect 433 1133 447 1147
rect 413 1113 427 1127
rect 433 1093 447 1107
rect 453 1093 467 1107
rect 393 1073 407 1087
rect 473 1073 487 1087
rect 353 1053 367 1067
rect 613 1553 627 1567
rect 653 1533 667 1547
rect 613 1313 627 1327
rect 653 1313 667 1327
rect 593 1273 607 1287
rect 613 1273 627 1287
rect 593 1253 607 1267
rect 573 1233 587 1247
rect 513 1213 527 1227
rect 573 1213 587 1227
rect 553 1193 567 1207
rect 533 1133 547 1147
rect 553 1133 567 1147
rect 633 1233 647 1247
rect 613 1193 627 1207
rect 593 1173 607 1187
rect 613 1173 627 1187
rect 653 1173 667 1187
rect 513 1093 527 1107
rect 553 1093 567 1107
rect 533 1073 547 1087
rect 573 1073 587 1087
rect 493 1053 507 1067
rect 533 1053 547 1067
rect 513 913 527 927
rect 493 893 507 907
rect 293 873 307 887
rect 413 873 427 887
rect 113 813 127 827
rect 133 813 147 827
rect 53 653 67 667
rect 253 853 267 867
rect 193 813 207 827
rect 153 793 167 807
rect 173 773 187 787
rect 233 813 247 827
rect 253 833 267 847
rect 373 853 387 867
rect 333 833 347 847
rect 213 693 227 707
rect 253 693 267 707
rect 153 673 167 687
rect 133 653 147 667
rect 193 653 207 667
rect 233 633 247 647
rect 133 613 147 627
rect 153 613 167 627
rect 193 613 207 627
rect 93 393 107 407
rect 173 593 187 607
rect 213 593 227 607
rect 233 413 247 427
rect 153 373 167 387
rect 93 333 107 347
rect 73 313 87 327
rect 33 193 47 207
rect 73 173 87 187
rect 193 373 207 387
rect 213 353 227 367
rect 353 813 367 827
rect 393 813 407 827
rect 293 773 307 787
rect 313 673 327 687
rect 353 673 367 687
rect 273 653 287 667
rect 273 633 287 647
rect 453 853 467 867
rect 433 793 447 807
rect 393 693 407 707
rect 413 693 427 707
rect 373 653 387 667
rect 353 633 367 647
rect 433 673 447 687
rect 313 613 327 627
rect 333 613 347 627
rect 293 593 307 607
rect 273 573 287 587
rect 393 613 407 627
rect 373 593 387 607
rect 313 513 327 527
rect 353 493 367 507
rect 313 453 327 467
rect 333 413 347 427
rect 253 353 267 367
rect 173 333 187 347
rect 293 333 307 347
rect 313 333 327 347
rect 253 313 267 327
rect 133 193 147 207
rect 233 193 247 207
rect 113 173 127 187
rect 93 153 107 167
rect 33 113 47 127
rect 73 133 87 147
rect 113 133 127 147
rect 153 133 167 147
rect 173 153 187 167
rect 393 433 407 447
rect 353 373 367 387
rect 373 373 387 387
rect 493 833 507 847
rect 493 793 507 807
rect 553 1033 567 1047
rect 573 893 587 907
rect 573 853 587 867
rect 593 833 607 847
rect 653 1153 667 1167
rect 713 1613 727 1627
rect 773 1633 787 1647
rect 693 1573 707 1587
rect 713 1573 727 1587
rect 693 1553 707 1567
rect 693 1493 707 1507
rect 733 1513 747 1527
rect 733 1453 747 1467
rect 713 1373 727 1387
rect 733 1333 747 1347
rect 713 1313 727 1327
rect 733 1293 747 1307
rect 713 1273 727 1287
rect 753 1273 767 1287
rect 693 1253 707 1267
rect 713 1213 727 1227
rect 713 1193 727 1207
rect 733 1173 747 1187
rect 813 1773 827 1787
rect 853 1773 867 1787
rect 873 1773 887 1787
rect 933 1773 947 1787
rect 813 1753 827 1767
rect 853 1753 867 1767
rect 873 1753 887 1767
rect 813 1713 827 1727
rect 853 1713 867 1727
rect 813 1613 827 1627
rect 793 1593 807 1607
rect 913 1733 927 1747
rect 1033 1853 1047 1867
rect 1013 1833 1027 1847
rect 1033 1833 1047 1847
rect 1073 1993 1087 2007
rect 993 1813 1007 1827
rect 973 1793 987 1807
rect 1033 1813 1047 1827
rect 1053 1813 1067 1827
rect 1193 2233 1207 2247
rect 1253 2213 1267 2227
rect 1213 2093 1227 2107
rect 1193 2053 1207 2067
rect 1213 2053 1227 2067
rect 1253 2073 1267 2087
rect 1453 2973 1467 2987
rect 1533 2973 1547 2987
rect 1453 2913 1467 2927
rect 1493 2913 1507 2927
rect 1573 2973 1587 2987
rect 1553 2853 1567 2867
rect 1453 2753 1467 2767
rect 1613 3033 1627 3047
rect 1593 2953 1607 2967
rect 1613 2953 1627 2967
rect 1573 2833 1587 2847
rect 1473 2673 1487 2687
rect 1433 2573 1447 2587
rect 1453 2573 1467 2587
rect 1493 2593 1507 2607
rect 1493 2573 1507 2587
rect 1433 2533 1447 2547
rect 1473 2553 1487 2567
rect 1393 2493 1407 2507
rect 1413 2493 1427 2507
rect 1353 2473 1367 2487
rect 1413 2473 1427 2487
rect 1313 2333 1327 2347
rect 1353 2333 1367 2347
rect 1313 2313 1327 2327
rect 1333 2233 1347 2247
rect 1313 2133 1327 2147
rect 1293 2073 1307 2087
rect 1273 2053 1287 2067
rect 1333 2073 1347 2087
rect 1313 2053 1327 2067
rect 1113 1993 1127 2007
rect 1173 1993 1187 2007
rect 1093 1833 1107 1847
rect 1093 1813 1107 1827
rect 1013 1773 1027 1787
rect 1033 1773 1047 1787
rect 953 1733 967 1747
rect 1013 1733 1027 1747
rect 1033 1733 1047 1747
rect 933 1693 947 1707
rect 973 1673 987 1687
rect 913 1633 927 1647
rect 913 1613 927 1627
rect 953 1613 967 1627
rect 873 1593 887 1607
rect 793 1573 807 1587
rect 813 1573 827 1587
rect 833 1573 847 1587
rect 813 1553 827 1567
rect 873 1573 887 1587
rect 913 1573 927 1587
rect 933 1573 947 1587
rect 853 1553 867 1567
rect 893 1553 907 1567
rect 793 1493 807 1507
rect 833 1473 847 1487
rect 813 1413 827 1427
rect 793 1333 807 1347
rect 793 1293 807 1307
rect 893 1513 907 1527
rect 913 1493 927 1507
rect 853 1453 867 1467
rect 873 1453 887 1467
rect 833 1353 847 1367
rect 833 1333 847 1347
rect 833 1293 847 1307
rect 813 1273 827 1287
rect 793 1213 807 1227
rect 793 1193 807 1207
rect 673 1073 687 1087
rect 633 1013 647 1027
rect 733 1113 747 1127
rect 733 1073 747 1087
rect 773 1113 787 1127
rect 773 1073 787 1087
rect 773 1013 787 1027
rect 773 993 787 1007
rect 753 913 767 927
rect 693 873 707 887
rect 653 853 667 867
rect 693 853 707 867
rect 733 853 747 867
rect 693 833 707 847
rect 633 793 647 807
rect 673 793 687 807
rect 713 793 727 807
rect 473 733 487 747
rect 533 733 547 747
rect 553 733 567 747
rect 533 713 547 727
rect 453 653 467 667
rect 433 493 447 507
rect 433 473 447 487
rect 493 633 507 647
rect 473 613 487 627
rect 493 593 507 607
rect 473 513 487 527
rect 433 393 447 407
rect 453 393 467 407
rect 513 573 527 587
rect 533 573 547 587
rect 593 753 607 767
rect 613 693 627 707
rect 573 633 587 647
rect 553 553 567 567
rect 513 493 527 507
rect 493 473 507 487
rect 513 453 527 467
rect 393 353 407 367
rect 413 333 427 347
rect 453 373 467 387
rect 493 373 507 387
rect 613 653 627 667
rect 653 753 667 767
rect 633 633 647 647
rect 693 773 707 787
rect 673 673 687 687
rect 753 813 767 827
rect 733 753 747 767
rect 633 613 647 627
rect 713 633 727 647
rect 613 493 627 507
rect 533 413 547 427
rect 593 413 607 427
rect 353 313 367 327
rect 433 313 447 327
rect 473 313 487 327
rect 513 313 527 327
rect 473 293 487 307
rect 353 273 367 287
rect 353 253 367 267
rect 253 173 267 187
rect 313 173 327 187
rect 333 173 347 187
rect 413 233 427 247
rect 273 133 287 147
rect 293 153 307 167
rect 313 153 327 167
rect 333 133 347 147
rect 373 153 387 167
rect 593 353 607 367
rect 553 253 567 267
rect 553 193 567 207
rect 433 173 447 187
rect 473 173 487 187
rect 533 173 547 187
rect 453 133 467 147
rect 493 153 507 167
rect 513 133 527 147
rect 693 533 707 547
rect 633 433 647 447
rect 653 393 667 407
rect 693 393 707 407
rect 713 333 727 347
rect 633 313 647 327
rect 693 313 707 327
rect 673 213 687 227
rect 613 193 627 207
rect 773 733 787 747
rect 853 1273 867 1287
rect 933 1413 947 1427
rect 953 1373 967 1387
rect 893 1353 907 1367
rect 853 1233 867 1247
rect 873 1233 887 1247
rect 853 1213 867 1227
rect 833 1153 847 1167
rect 833 1133 847 1147
rect 813 1113 827 1127
rect 993 1633 1007 1647
rect 1013 1593 1027 1607
rect 1073 1753 1087 1767
rect 1153 1853 1167 1867
rect 1153 1813 1167 1827
rect 1133 1773 1147 1787
rect 1013 1573 1027 1587
rect 1013 1553 1027 1567
rect 1053 1553 1067 1567
rect 993 1533 1007 1547
rect 1033 1533 1047 1547
rect 1173 1733 1187 1747
rect 1133 1653 1147 1667
rect 1113 1633 1127 1647
rect 1113 1573 1127 1587
rect 1153 1573 1167 1587
rect 1173 1593 1187 1607
rect 1193 1593 1207 1607
rect 1293 2013 1307 2027
rect 1233 1833 1247 1847
rect 1273 1833 1287 1847
rect 1293 1833 1307 1847
rect 1253 1813 1267 1827
rect 1233 1753 1247 1767
rect 1293 1813 1307 1827
rect 1293 1773 1307 1787
rect 1273 1733 1287 1747
rect 1253 1713 1267 1727
rect 1273 1693 1287 1707
rect 1253 1673 1267 1687
rect 1213 1573 1227 1587
rect 1233 1573 1247 1587
rect 1093 1553 1107 1567
rect 1153 1553 1167 1567
rect 1173 1553 1187 1567
rect 1213 1553 1227 1567
rect 1433 2413 1447 2427
rect 1513 2513 1527 2527
rect 1533 2533 1547 2547
rect 1553 2513 1567 2527
rect 1493 2373 1507 2387
rect 1473 2353 1487 2367
rect 1473 2333 1487 2347
rect 1413 2253 1427 2267
rect 1373 2193 1387 2207
rect 1453 2253 1467 2267
rect 1613 2813 1627 2827
rect 1693 3213 1707 3227
rect 1713 3213 1727 3227
rect 1713 3193 1727 3207
rect 1693 3153 1707 3167
rect 1653 3093 1667 3107
rect 1733 3133 1747 3147
rect 1733 3113 1747 3127
rect 1713 3073 1727 3087
rect 1653 2973 1667 2987
rect 1633 2773 1647 2787
rect 1633 2693 1647 2707
rect 1693 2993 1707 3007
rect 1813 3453 1827 3467
rect 1853 3433 1867 3447
rect 1773 3393 1787 3407
rect 1793 3373 1807 3387
rect 1833 3293 1847 3307
rect 1813 3273 1827 3287
rect 1913 3633 1927 3647
rect 1933 3613 1947 3627
rect 1893 3473 1907 3487
rect 1913 3473 1927 3487
rect 1893 3433 1907 3447
rect 1833 3253 1847 3267
rect 1793 3213 1807 3227
rect 1893 3253 1907 3267
rect 1833 3213 1847 3227
rect 1873 3213 1887 3227
rect 1893 3213 1907 3227
rect 1833 3193 1847 3207
rect 1873 3193 1887 3207
rect 1773 3153 1787 3167
rect 1793 3153 1807 3167
rect 1753 3093 1767 3107
rect 1813 3133 1827 3147
rect 1753 3033 1767 3047
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1793 2993 1807 3007
rect 1993 3593 2007 3607
rect 2293 3973 2307 3987
rect 2153 3733 2167 3747
rect 1953 3473 1967 3487
rect 1973 3473 1987 3487
rect 1993 3493 2007 3507
rect 2013 3453 2027 3467
rect 1973 3373 1987 3387
rect 1933 3353 1947 3367
rect 1953 3273 1967 3287
rect 1973 3253 1987 3267
rect 1933 3213 1947 3227
rect 1913 3133 1927 3147
rect 1853 3093 1867 3107
rect 1873 3093 1887 3107
rect 1893 3033 1907 3047
rect 1873 3013 1887 3027
rect 1833 2993 1847 3007
rect 1693 2913 1707 2927
rect 1693 2893 1707 2907
rect 1673 2873 1687 2887
rect 1693 2813 1707 2827
rect 1693 2673 1707 2687
rect 1653 2653 1667 2667
rect 1673 2633 1687 2647
rect 1653 2613 1667 2627
rect 1593 2593 1607 2607
rect 1593 2513 1607 2527
rect 1593 2493 1607 2507
rect 1573 2333 1587 2347
rect 1553 2273 1567 2287
rect 1573 2253 1587 2267
rect 1573 2233 1587 2247
rect 1413 2093 1427 2107
rect 1373 2073 1387 2087
rect 1353 1973 1367 1987
rect 1433 2033 1447 2047
rect 1393 2013 1407 2027
rect 1533 2213 1547 2227
rect 1553 2073 1567 2087
rect 1493 2053 1507 2067
rect 1533 2033 1547 2047
rect 1513 1993 1527 2007
rect 1573 1993 1587 2007
rect 1393 1913 1407 1927
rect 1453 1913 1467 1927
rect 1313 1693 1327 1707
rect 1293 1673 1307 1687
rect 1373 1713 1387 1727
rect 1353 1653 1367 1667
rect 1313 1613 1327 1627
rect 1333 1613 1347 1627
rect 1373 1613 1387 1627
rect 1273 1553 1287 1567
rect 993 1493 1007 1507
rect 1033 1433 1047 1447
rect 973 1353 987 1367
rect 913 1333 927 1347
rect 933 1313 947 1327
rect 973 1333 987 1347
rect 1013 1333 1027 1347
rect 1033 1333 1047 1347
rect 913 1293 927 1307
rect 913 1273 927 1287
rect 993 1273 1007 1287
rect 893 1213 907 1227
rect 893 1153 907 1167
rect 853 1093 867 1107
rect 993 1253 1007 1267
rect 993 1193 1007 1207
rect 973 1153 987 1167
rect 1093 1353 1107 1367
rect 1073 1333 1087 1347
rect 1113 1333 1127 1347
rect 1093 1313 1107 1327
rect 1113 1313 1127 1327
rect 1093 1293 1107 1307
rect 1053 1253 1067 1267
rect 1053 1193 1067 1207
rect 1033 1173 1047 1187
rect 1033 1133 1047 1147
rect 933 1113 947 1127
rect 1093 1153 1107 1167
rect 1053 1093 1067 1107
rect 953 1073 967 1087
rect 873 1053 887 1067
rect 893 1053 907 1067
rect 813 1013 827 1027
rect 833 973 847 987
rect 813 913 827 927
rect 853 893 867 907
rect 833 853 847 867
rect 833 813 847 827
rect 853 813 867 827
rect 813 693 827 707
rect 793 673 807 687
rect 833 653 847 667
rect 813 633 827 647
rect 773 593 787 607
rect 773 533 787 547
rect 893 973 907 987
rect 993 953 1007 967
rect 893 933 907 947
rect 913 893 927 907
rect 893 853 907 867
rect 953 853 967 867
rect 973 853 987 867
rect 893 813 907 827
rect 973 813 987 827
rect 933 793 947 807
rect 873 773 887 787
rect 1073 953 1087 967
rect 1073 933 1087 947
rect 1013 913 1027 927
rect 1073 873 1087 887
rect 1193 1533 1207 1547
rect 1233 1533 1247 1547
rect 1253 1533 1267 1547
rect 1293 1513 1307 1527
rect 1333 1573 1347 1587
rect 1333 1553 1347 1567
rect 1233 1493 1247 1507
rect 1313 1493 1327 1507
rect 1193 1473 1207 1487
rect 1173 1433 1187 1447
rect 1253 1393 1267 1407
rect 1193 1373 1207 1387
rect 1173 1333 1187 1347
rect 1213 1353 1227 1367
rect 1193 1313 1207 1327
rect 1153 1293 1167 1307
rect 1193 1233 1207 1247
rect 1193 1213 1207 1227
rect 1133 1193 1147 1207
rect 1273 1333 1287 1347
rect 1253 1293 1267 1307
rect 1173 1173 1187 1187
rect 1213 1173 1227 1187
rect 1133 1153 1147 1167
rect 1113 1133 1127 1147
rect 1193 1153 1207 1167
rect 1113 1113 1127 1127
rect 1153 1073 1167 1087
rect 1153 973 1167 987
rect 1173 953 1187 967
rect 1113 913 1127 927
rect 1013 853 1027 867
rect 1053 853 1067 867
rect 1093 853 1107 867
rect 1113 853 1127 867
rect 1053 833 1067 847
rect 1033 753 1047 767
rect 993 713 1007 727
rect 893 693 907 707
rect 953 693 967 707
rect 873 653 887 667
rect 853 633 867 647
rect 913 673 927 687
rect 1013 673 1027 687
rect 993 653 1007 667
rect 893 613 907 627
rect 933 613 947 627
rect 973 613 987 627
rect 853 593 867 607
rect 873 593 887 607
rect 893 573 907 587
rect 873 453 887 467
rect 873 413 887 427
rect 773 353 787 367
rect 853 393 867 407
rect 973 433 987 447
rect 933 393 947 407
rect 833 373 847 387
rect 893 373 907 387
rect 953 353 967 367
rect 813 333 827 347
rect 793 313 807 327
rect 753 293 767 307
rect 733 233 747 247
rect 813 293 827 307
rect 913 313 927 327
rect 953 273 967 287
rect 913 253 927 267
rect 893 233 907 247
rect 813 213 827 227
rect 853 213 867 227
rect 893 213 907 227
rect 633 173 647 187
rect 593 153 607 167
rect 553 133 567 147
rect 853 193 867 207
rect 753 173 767 187
rect 773 173 787 187
rect 793 173 807 187
rect 733 153 747 167
rect 753 133 767 147
rect 793 133 807 147
rect 833 133 847 147
rect 593 113 607 127
rect 653 113 667 127
rect 613 93 627 107
rect 833 93 847 107
rect 873 153 887 167
rect 1093 813 1107 827
rect 1253 1253 1267 1267
rect 1233 1133 1247 1147
rect 1213 1073 1227 1087
rect 1233 1093 1247 1107
rect 1253 953 1267 967
rect 1193 933 1207 947
rect 1193 913 1207 927
rect 1213 893 1227 907
rect 1433 1873 1447 1887
rect 1433 1813 1447 1827
rect 1533 1813 1547 1827
rect 1413 1773 1427 1787
rect 1473 1793 1487 1807
rect 1533 1793 1547 1807
rect 1553 1793 1567 1807
rect 1513 1773 1527 1787
rect 1493 1753 1507 1767
rect 1453 1733 1467 1747
rect 1473 1633 1487 1647
rect 1533 1633 1547 1647
rect 1573 1633 1587 1647
rect 1413 1573 1427 1587
rect 1413 1553 1427 1567
rect 1633 2533 1647 2547
rect 1653 2513 1667 2527
rect 1633 2373 1647 2387
rect 1613 2273 1627 2287
rect 1693 2553 1707 2567
rect 1673 2473 1687 2487
rect 1793 2933 1807 2947
rect 1753 2873 1767 2887
rect 1753 2793 1767 2807
rect 1773 2793 1787 2807
rect 1753 2733 1767 2747
rect 1833 2773 1847 2787
rect 1813 2753 1827 2767
rect 1853 2753 1867 2767
rect 1833 2733 1847 2747
rect 1853 2733 1867 2747
rect 1773 2673 1787 2687
rect 1853 2693 1867 2707
rect 1833 2653 1847 2667
rect 1733 2553 1747 2567
rect 1653 2253 1667 2267
rect 1673 2213 1687 2227
rect 1793 2593 1807 2607
rect 1813 2513 1827 2527
rect 1813 2493 1827 2507
rect 1793 2473 1807 2487
rect 1853 2473 1867 2487
rect 1993 3173 2007 3187
rect 2033 3273 2047 3287
rect 2133 3693 2147 3707
rect 2333 3733 2347 3747
rect 2153 3593 2167 3607
rect 2313 3713 2327 3727
rect 2313 3593 2327 3607
rect 2173 3573 2187 3587
rect 2173 3553 2187 3567
rect 2293 3553 2307 3567
rect 2113 3533 2127 3547
rect 2113 3513 2127 3527
rect 2153 3513 2167 3527
rect 2233 3513 2247 3527
rect 2113 3473 2127 3487
rect 2253 3493 2267 3507
rect 2093 3453 2107 3467
rect 2093 3413 2107 3427
rect 2073 3253 2087 3267
rect 2153 3333 2167 3347
rect 2133 3313 2147 3327
rect 2113 3253 2127 3267
rect 2033 3213 2047 3227
rect 2073 3213 2087 3227
rect 2133 3233 2147 3247
rect 2153 3233 2167 3247
rect 2113 3213 2127 3227
rect 1973 3133 1987 3147
rect 1953 3113 1967 3127
rect 1933 3053 1947 3067
rect 2073 3193 2087 3207
rect 1913 2833 1927 2847
rect 1893 2793 1907 2807
rect 1973 2993 1987 3007
rect 2033 3093 2047 3107
rect 2093 3073 2107 3087
rect 2153 3113 2167 3127
rect 2133 3073 2147 3087
rect 2113 3053 2127 3067
rect 2053 3013 2067 3027
rect 2073 3013 2087 3027
rect 2113 3013 2127 3027
rect 2133 3033 2147 3047
rect 2273 3293 2287 3307
rect 2273 3273 2287 3287
rect 2193 3213 2207 3227
rect 2213 3233 2227 3247
rect 2253 3233 2267 3247
rect 2333 3493 2347 3507
rect 2373 3913 2387 3927
rect 2373 3693 2387 3707
rect 2393 3653 2407 3667
rect 2373 3613 2387 3627
rect 2373 3533 2387 3547
rect 2613 3973 2627 3987
rect 2473 3893 2487 3907
rect 2473 3733 2487 3747
rect 2493 3693 2507 3707
rect 2533 3693 2547 3707
rect 2453 3673 2467 3687
rect 2493 3573 2507 3587
rect 2433 3553 2447 3567
rect 2393 3493 2407 3507
rect 2353 3353 2367 3367
rect 2333 3293 2347 3307
rect 2393 3293 2407 3307
rect 2293 3253 2307 3267
rect 2353 3273 2367 3287
rect 2233 3213 2247 3227
rect 2273 3213 2287 3227
rect 2173 3093 2187 3107
rect 2273 3073 2287 3087
rect 2193 3033 2207 3047
rect 2153 3013 2167 3027
rect 2233 3033 2247 3047
rect 2213 3013 2227 3027
rect 2073 2993 2087 3007
rect 2013 2953 2027 2967
rect 2013 2793 2027 2807
rect 2053 2793 2067 2807
rect 1973 2773 1987 2787
rect 1893 2753 1907 2767
rect 1933 2753 1947 2767
rect 1993 2733 2007 2747
rect 1893 2713 1907 2727
rect 1913 2673 1927 2687
rect 1953 2693 1967 2707
rect 1933 2553 1947 2567
rect 1893 2493 1907 2507
rect 1773 2413 1787 2427
rect 1813 2453 1827 2467
rect 1793 2253 1807 2267
rect 1833 2233 1847 2247
rect 1873 2213 1887 2227
rect 1713 2193 1727 2207
rect 1813 2193 1827 2207
rect 1633 2173 1647 2187
rect 1693 2173 1707 2187
rect 1773 2173 1787 2187
rect 1693 2153 1707 2167
rect 1653 2113 1667 2127
rect 1753 2133 1767 2147
rect 1733 2093 1747 2107
rect 1753 2093 1767 2107
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1693 2073 1707 2087
rect 1813 2153 1827 2167
rect 1833 2153 1847 2167
rect 1873 2153 1887 2167
rect 1853 2093 1867 2107
rect 1713 2053 1727 2067
rect 1733 2053 1747 2067
rect 1753 2053 1767 2067
rect 1653 1973 1667 1987
rect 1613 1813 1627 1827
rect 1633 1793 1647 1807
rect 1633 1753 1647 1767
rect 1613 1673 1627 1687
rect 1533 1613 1547 1627
rect 1593 1613 1607 1627
rect 1493 1573 1507 1587
rect 1513 1553 1527 1567
rect 1433 1493 1447 1507
rect 1453 1493 1467 1507
rect 1413 1473 1427 1487
rect 1433 1413 1447 1427
rect 1393 1393 1407 1407
rect 1413 1393 1427 1407
rect 1373 1353 1387 1367
rect 1393 1353 1407 1367
rect 1293 1293 1307 1307
rect 1333 1313 1347 1327
rect 1313 1273 1327 1287
rect 1333 1253 1347 1267
rect 1293 1133 1307 1147
rect 1293 1113 1307 1127
rect 1313 1053 1327 1067
rect 1293 1013 1307 1027
rect 1213 873 1227 887
rect 1273 873 1287 887
rect 1193 833 1207 847
rect 1313 913 1327 927
rect 1373 1253 1387 1267
rect 1353 1193 1367 1207
rect 1353 1133 1367 1147
rect 1393 1213 1407 1227
rect 1373 1113 1387 1127
rect 1493 1473 1507 1487
rect 1473 1373 1487 1387
rect 1453 1333 1467 1347
rect 1513 1433 1527 1447
rect 1493 1353 1507 1367
rect 1553 1573 1567 1587
rect 1573 1573 1587 1587
rect 1613 1593 1627 1607
rect 1733 2013 1747 2027
rect 2053 2693 2067 2707
rect 2033 2673 2047 2687
rect 2253 2833 2267 2847
rect 2233 2793 2247 2807
rect 2213 2773 2227 2787
rect 2153 2753 2167 2767
rect 2133 2733 2147 2747
rect 2333 3233 2347 3247
rect 2333 3193 2347 3207
rect 2393 3213 2407 3227
rect 2373 3133 2387 3147
rect 2353 3093 2367 3107
rect 2293 3033 2307 3047
rect 2353 3033 2367 3047
rect 2293 2993 2307 3007
rect 2313 3013 2327 3027
rect 2373 3013 2387 3027
rect 2433 3533 2447 3547
rect 2453 3213 2467 3227
rect 2453 3173 2467 3187
rect 2453 3073 2467 3087
rect 2433 3053 2447 3067
rect 2413 3013 2427 3027
rect 2333 2993 2347 3007
rect 2393 2993 2407 3007
rect 2353 2773 2367 2787
rect 2093 2713 2107 2727
rect 2273 2753 2287 2767
rect 2333 2753 2347 2767
rect 2193 2713 2207 2727
rect 2253 2713 2267 2727
rect 2273 2693 2287 2707
rect 2313 2713 2327 2727
rect 2093 2673 2107 2687
rect 2113 2673 2127 2687
rect 2293 2673 2307 2687
rect 2073 2633 2087 2647
rect 2273 2653 2287 2667
rect 2193 2633 2207 2647
rect 1973 2573 1987 2587
rect 2073 2573 2087 2587
rect 2133 2573 2147 2587
rect 2013 2533 2027 2547
rect 1993 2513 2007 2527
rect 2113 2553 2127 2567
rect 2093 2533 2107 2547
rect 2053 2513 2067 2527
rect 2033 2493 2047 2507
rect 1953 2473 1967 2487
rect 2033 2473 2047 2487
rect 1933 2413 1947 2427
rect 1973 2293 1987 2307
rect 1913 2273 1927 2287
rect 1973 2273 1987 2287
rect 2013 2273 2027 2287
rect 1913 2233 1927 2247
rect 1953 2213 1967 2227
rect 1933 2193 1947 2207
rect 1933 2153 1947 2167
rect 1893 2113 1907 2127
rect 1913 2113 1927 2127
rect 1993 2173 2007 2187
rect 1973 2113 1987 2127
rect 1933 2093 1947 2107
rect 1953 2093 1967 2107
rect 2253 2573 2267 2587
rect 2293 2633 2307 2647
rect 2173 2533 2187 2547
rect 2193 2533 2207 2547
rect 2213 2533 2227 2547
rect 2093 2453 2107 2467
rect 2073 2293 2087 2307
rect 2053 2133 2067 2147
rect 2053 2113 2067 2127
rect 1913 2073 1927 2087
rect 1953 2053 1967 2067
rect 2033 2073 2047 2087
rect 2153 2413 2167 2427
rect 2113 2213 2127 2227
rect 2253 2353 2267 2367
rect 2213 2273 2227 2287
rect 2193 2213 2207 2227
rect 2173 2173 2187 2187
rect 2153 2133 2167 2147
rect 2113 2073 2127 2087
rect 1933 2033 1947 2047
rect 1893 2013 1907 2027
rect 1873 1993 1887 2007
rect 1713 1893 1727 1907
rect 1753 1893 1767 1907
rect 1713 1833 1727 1847
rect 1673 1813 1687 1827
rect 1653 1733 1667 1747
rect 1913 1973 1927 1987
rect 1713 1793 1727 1807
rect 1793 1813 1807 1827
rect 1793 1793 1807 1807
rect 1733 1773 1747 1787
rect 1693 1693 1707 1707
rect 1673 1613 1687 1627
rect 1553 1453 1567 1467
rect 1533 1413 1547 1427
rect 1553 1393 1567 1407
rect 1513 1333 1527 1347
rect 1433 1313 1447 1327
rect 1453 1293 1467 1307
rect 1533 1313 1547 1327
rect 1493 1273 1507 1287
rect 1533 1253 1547 1267
rect 1553 1253 1567 1267
rect 1413 1113 1427 1127
rect 1433 1113 1447 1127
rect 1353 1073 1367 1087
rect 1373 1073 1387 1087
rect 1413 1073 1427 1087
rect 1353 913 1367 927
rect 1393 1053 1407 1067
rect 1513 1153 1527 1167
rect 1473 1113 1487 1127
rect 1493 1093 1507 1107
rect 1453 1073 1467 1087
rect 1473 1073 1487 1087
rect 1433 973 1447 987
rect 1433 913 1447 927
rect 1393 893 1407 907
rect 1373 873 1387 887
rect 1333 853 1347 867
rect 1373 853 1387 867
rect 1253 833 1267 847
rect 1293 833 1307 847
rect 1333 833 1347 847
rect 1093 793 1107 807
rect 1073 773 1087 787
rect 1033 653 1047 667
rect 1053 653 1067 667
rect 1013 633 1027 647
rect 1133 753 1147 767
rect 1293 773 1307 787
rect 1273 753 1287 767
rect 1233 733 1247 747
rect 1233 713 1247 727
rect 1413 833 1427 847
rect 1353 793 1367 807
rect 1393 753 1407 767
rect 1413 753 1427 767
rect 1193 693 1207 707
rect 1113 673 1127 687
rect 1053 633 1067 647
rect 1013 613 1027 627
rect 1073 613 1087 627
rect 1093 633 1107 647
rect 1133 633 1147 647
rect 1113 613 1127 627
rect 1313 693 1327 707
rect 1333 693 1347 707
rect 1273 673 1287 687
rect 1173 613 1187 627
rect 1213 613 1227 627
rect 1253 613 1267 627
rect 1073 593 1087 607
rect 993 413 1007 427
rect 1113 533 1127 547
rect 1153 533 1167 547
rect 1073 493 1087 507
rect 1213 493 1227 507
rect 1133 413 1147 427
rect 1013 353 1027 367
rect 1113 373 1127 387
rect 1173 393 1187 407
rect 1353 673 1367 687
rect 1453 893 1467 907
rect 1433 733 1447 747
rect 1433 673 1447 687
rect 1673 1573 1687 1587
rect 1693 1573 1707 1587
rect 1633 1553 1647 1567
rect 1773 1753 1787 1767
rect 1813 1773 1827 1787
rect 1853 1773 1867 1787
rect 1993 2013 2007 2027
rect 1933 1813 1947 1827
rect 1833 1753 1847 1767
rect 1833 1713 1847 1727
rect 1853 1653 1867 1667
rect 1833 1613 1847 1627
rect 1753 1593 1767 1607
rect 1813 1593 1827 1607
rect 1833 1593 1847 1607
rect 1753 1553 1767 1567
rect 1613 1513 1627 1527
rect 1593 1493 1607 1507
rect 1693 1473 1707 1487
rect 1673 1353 1687 1367
rect 1593 1293 1607 1307
rect 1613 1313 1627 1327
rect 1573 1233 1587 1247
rect 1573 1173 1587 1187
rect 1553 1113 1567 1127
rect 1553 1093 1567 1107
rect 1573 1033 1587 1047
rect 1533 993 1547 1007
rect 1493 973 1507 987
rect 1533 933 1547 947
rect 1613 1193 1627 1207
rect 1653 1273 1667 1287
rect 1633 1173 1647 1187
rect 1733 1393 1747 1407
rect 1793 1553 1807 1567
rect 1833 1553 1847 1567
rect 1773 1533 1787 1547
rect 1793 1473 1807 1487
rect 1953 1633 1967 1647
rect 1913 1613 1927 1627
rect 1933 1613 1947 1627
rect 1873 1593 1887 1607
rect 1913 1573 1927 1587
rect 1953 1573 1967 1587
rect 1893 1553 1907 1567
rect 1853 1533 1867 1547
rect 1833 1393 1847 1407
rect 1853 1393 1867 1407
rect 1753 1333 1767 1347
rect 1773 1313 1787 1327
rect 1693 1293 1707 1307
rect 1813 1313 1827 1327
rect 1713 1273 1727 1287
rect 1793 1273 1807 1287
rect 1693 1253 1707 1267
rect 1773 1193 1787 1207
rect 1693 1153 1707 1167
rect 1613 1133 1627 1147
rect 1633 1133 1647 1147
rect 1673 1133 1687 1147
rect 1693 1133 1707 1147
rect 1673 1113 1687 1127
rect 1613 1073 1627 1087
rect 1653 1073 1667 1087
rect 1753 1113 1767 1127
rect 1713 1093 1727 1107
rect 1733 1073 1747 1087
rect 1613 1053 1627 1067
rect 1633 1013 1647 1027
rect 1613 913 1627 927
rect 1553 873 1567 887
rect 1593 873 1607 887
rect 1473 853 1487 867
rect 1533 853 1547 867
rect 1553 833 1567 847
rect 1573 853 1587 867
rect 1553 813 1567 827
rect 1593 813 1607 827
rect 1493 773 1507 787
rect 1473 733 1487 747
rect 1453 653 1467 667
rect 1493 693 1507 707
rect 1293 613 1307 627
rect 1373 633 1387 647
rect 1413 633 1427 647
rect 1373 593 1387 607
rect 1353 513 1367 527
rect 1273 433 1287 447
rect 1353 433 1367 447
rect 1533 673 1547 687
rect 1513 653 1527 667
rect 1453 593 1467 607
rect 1413 573 1427 587
rect 1493 533 1507 547
rect 1513 533 1527 547
rect 1753 1033 1767 1047
rect 1653 993 1667 1007
rect 1753 973 1767 987
rect 1653 933 1667 947
rect 1633 893 1647 907
rect 1653 893 1667 907
rect 1733 873 1747 887
rect 1673 833 1687 847
rect 1713 813 1727 827
rect 1613 753 1627 767
rect 1713 793 1727 807
rect 1713 773 1727 787
rect 1693 713 1707 727
rect 1653 693 1667 707
rect 1833 1253 1847 1267
rect 1933 1373 1947 1387
rect 1913 1353 1927 1367
rect 1873 1293 1887 1307
rect 1853 1213 1867 1227
rect 1793 1133 1807 1147
rect 1853 1133 1867 1147
rect 1913 1313 1927 1327
rect 1933 1333 1947 1347
rect 1893 1273 1907 1287
rect 1873 1113 1887 1127
rect 1933 1293 1947 1307
rect 2013 1993 2027 2007
rect 2093 2053 2107 2067
rect 2273 2313 2287 2327
rect 2253 2273 2267 2287
rect 2253 2253 2267 2267
rect 2333 2573 2347 2587
rect 2313 2533 2327 2547
rect 2333 2513 2347 2527
rect 2453 3013 2467 3027
rect 2473 3013 2487 3027
rect 2453 2973 2467 2987
rect 2753 4113 2767 4127
rect 3013 4513 3027 4527
rect 3053 4513 3067 4527
rect 3093 4513 3107 4527
rect 2933 4493 2947 4507
rect 2993 4493 3007 4507
rect 2973 4453 2987 4467
rect 3173 4513 3187 4527
rect 3233 4513 3247 4527
rect 3113 4493 3127 4507
rect 3133 4493 3147 4507
rect 3173 4493 3187 4507
rect 3033 4453 3047 4467
rect 3073 4453 3087 4467
rect 3113 4453 3127 4467
rect 3073 4433 3087 4447
rect 3013 4413 3027 4427
rect 2913 4213 2927 4227
rect 2873 4193 2887 4207
rect 2853 4153 2867 4167
rect 2933 4173 2947 4187
rect 2973 4173 2987 4187
rect 3013 4193 3027 4207
rect 3053 4193 3067 4207
rect 2953 4153 2967 4167
rect 2913 4133 2927 4147
rect 2953 4133 2967 4147
rect 2993 4133 3007 4147
rect 2713 4073 2727 4087
rect 2813 4073 2827 4087
rect 2673 3953 2687 3967
rect 2733 4033 2747 4047
rect 2773 3993 2787 4007
rect 2773 3953 2787 3967
rect 3253 4453 3267 4467
rect 3273 4473 3287 4487
rect 3413 4493 3427 4507
rect 3293 4453 3307 4467
rect 3353 4473 3367 4487
rect 3373 4473 3387 4487
rect 3393 4453 3407 4467
rect 3193 4413 3207 4427
rect 3193 4273 3207 4287
rect 3113 4253 3127 4267
rect 3253 4253 3267 4267
rect 3093 4213 3107 4227
rect 3113 4193 3127 4207
rect 3073 4153 3087 4167
rect 3093 4153 3107 4167
rect 3033 4113 3047 4127
rect 2993 4033 3007 4047
rect 3053 4013 3067 4027
rect 3073 4013 3087 4027
rect 2633 3713 2647 3727
rect 2613 3693 2627 3707
rect 2673 3713 2687 3727
rect 2713 3693 2727 3707
rect 2653 3673 2667 3687
rect 2673 3673 2687 3687
rect 2753 3673 2767 3687
rect 2593 3653 2607 3667
rect 2573 3553 2587 3567
rect 2533 3533 2547 3547
rect 2513 3353 2527 3367
rect 2753 3653 2767 3667
rect 2913 3973 2927 3987
rect 2973 3973 2987 3987
rect 3233 4213 3247 4227
rect 3213 4173 3227 4187
rect 3273 4233 3287 4247
rect 3393 4233 3407 4247
rect 3293 4193 3307 4207
rect 3313 4213 3327 4227
rect 3253 4153 3267 4167
rect 3333 4153 3347 4167
rect 3373 4153 3387 4167
rect 3153 4113 3167 4127
rect 3353 4053 3367 4067
rect 3233 4033 3247 4047
rect 3213 4013 3227 4027
rect 3013 3973 3027 3987
rect 3093 3993 3107 4007
rect 2933 3953 2947 3967
rect 2873 3693 2887 3707
rect 2793 3673 2807 3687
rect 2913 3693 2927 3707
rect 2893 3673 2907 3687
rect 2813 3633 2827 3647
rect 2773 3613 2787 3627
rect 2913 3613 2927 3627
rect 2713 3553 2727 3567
rect 2673 3513 2687 3527
rect 2693 3493 2707 3507
rect 2733 3493 2747 3507
rect 2553 3193 2567 3207
rect 2513 3113 2527 3127
rect 2513 3033 2527 3047
rect 2673 3153 2687 3167
rect 2633 3133 2647 3147
rect 2613 3053 2627 3067
rect 2533 3013 2547 3027
rect 2533 2993 2547 3007
rect 2493 2813 2507 2827
rect 2473 2793 2487 2807
rect 2493 2793 2507 2807
rect 2433 2773 2447 2787
rect 2473 2773 2487 2787
rect 2373 2753 2387 2767
rect 2413 2753 2427 2767
rect 2433 2733 2447 2747
rect 2393 2633 2407 2647
rect 2373 2593 2387 2607
rect 2453 2693 2467 2707
rect 2473 2573 2487 2587
rect 2513 2733 2527 2747
rect 2593 2973 2607 2987
rect 2813 3513 2827 3527
rect 2833 3513 2847 3527
rect 2873 3493 2887 3507
rect 2893 3473 2907 3487
rect 2753 3413 2767 3427
rect 2713 3173 2727 3187
rect 2713 3093 2727 3107
rect 2773 3213 2787 3227
rect 2833 3213 2847 3227
rect 2773 3153 2787 3167
rect 2753 3053 2767 3067
rect 2653 3033 2667 3047
rect 2673 3033 2687 3047
rect 2693 3033 2707 3047
rect 2713 3013 2727 3027
rect 2733 2993 2747 3007
rect 2633 2793 2647 2807
rect 2553 2773 2567 2787
rect 2593 2773 2607 2787
rect 2553 2733 2567 2747
rect 2573 2733 2587 2747
rect 2633 2753 2647 2767
rect 2793 3053 2807 3067
rect 2773 2853 2787 2867
rect 2733 2753 2747 2767
rect 2773 2753 2787 2767
rect 2753 2733 2767 2747
rect 2533 2693 2547 2707
rect 2513 2653 2527 2667
rect 2393 2553 2407 2567
rect 2373 2533 2387 2547
rect 2413 2533 2427 2547
rect 2493 2553 2507 2567
rect 2653 2713 2667 2727
rect 2713 2713 2727 2727
rect 2853 3193 2867 3207
rect 2893 3153 2907 3167
rect 2853 3093 2867 3107
rect 2873 3093 2887 3107
rect 2893 3093 2907 3107
rect 2853 3073 2867 3087
rect 2833 2993 2847 3007
rect 2813 2793 2827 2807
rect 2833 2753 2847 2767
rect 2853 2773 2867 2787
rect 3133 3953 3147 3967
rect 3153 3973 3167 3987
rect 3173 3933 3187 3947
rect 3153 3753 3167 3767
rect 3273 4013 3287 4027
rect 3313 4013 3327 4027
rect 3333 4013 3347 4027
rect 3253 3973 3267 3987
rect 2973 3713 2987 3727
rect 2953 3673 2967 3687
rect 2953 3653 2967 3667
rect 2993 3633 3007 3647
rect 3153 3713 3167 3727
rect 3213 3713 3227 3727
rect 3073 3673 3087 3687
rect 3113 3653 3127 3667
rect 3133 3633 3147 3647
rect 3053 3593 3067 3607
rect 3193 3673 3207 3687
rect 3173 3573 3187 3587
rect 2933 3513 2947 3527
rect 2953 3473 2967 3487
rect 3033 3533 3047 3547
rect 3073 3513 3087 3527
rect 2993 3453 3007 3467
rect 2953 3233 2967 3247
rect 2973 3213 2987 3227
rect 2973 3113 2987 3127
rect 3213 3553 3227 3567
rect 3273 3733 3287 3747
rect 3353 3993 3367 4007
rect 3373 3993 3387 4007
rect 3353 3953 3367 3967
rect 3373 3953 3387 3967
rect 3453 4473 3467 4487
rect 3493 4513 3507 4527
rect 3433 4153 3447 4167
rect 3493 4233 3507 4247
rect 3493 4173 3507 4187
rect 3573 4473 3587 4487
rect 3633 4493 3647 4507
rect 3613 4213 3627 4227
rect 3613 4173 3627 4187
rect 3553 4093 3567 4107
rect 3533 4073 3547 4087
rect 3453 4013 3467 4027
rect 3473 4013 3487 4027
rect 3413 3993 3427 4007
rect 3433 3993 3447 4007
rect 3393 3733 3407 3747
rect 3253 3693 3267 3707
rect 3273 3713 3287 3727
rect 3293 3713 3307 3727
rect 3313 3713 3327 3727
rect 3333 3713 3347 3727
rect 3373 3673 3387 3687
rect 3353 3653 3367 3667
rect 3293 3613 3307 3627
rect 3273 3553 3287 3567
rect 3353 3553 3367 3567
rect 3153 3533 3167 3547
rect 3213 3533 3227 3547
rect 3233 3533 3247 3547
rect 3133 3513 3147 3527
rect 3093 3273 3107 3287
rect 3173 3513 3187 3527
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3253 3513 3267 3527
rect 3173 3473 3187 3487
rect 3233 3453 3247 3467
rect 3153 3313 3167 3327
rect 3313 3533 3327 3547
rect 3333 3533 3347 3547
rect 3393 3633 3407 3647
rect 3513 3973 3527 3987
rect 3573 3933 3587 3947
rect 3693 4453 3707 4467
rect 3713 4473 3727 4487
rect 3733 4453 3747 4467
rect 3653 4433 3667 4447
rect 3773 4433 3787 4447
rect 3793 4453 3807 4467
rect 3793 4413 3807 4427
rect 3653 4233 3667 4247
rect 3713 4233 3727 4247
rect 3673 4213 3687 4227
rect 3653 4153 3667 4167
rect 3773 4173 3787 4187
rect 3733 4153 3747 4167
rect 3773 4153 3787 4167
rect 3693 4093 3707 4107
rect 3653 4073 3667 4087
rect 3673 4033 3687 4047
rect 3693 3993 3707 4007
rect 3673 3953 3687 3967
rect 3633 3913 3647 3927
rect 3753 4013 3767 4027
rect 3773 3893 3787 3907
rect 3673 3833 3687 3847
rect 3513 3753 3527 3767
rect 3613 3753 3627 3767
rect 3433 3673 3447 3687
rect 3453 3653 3467 3667
rect 3413 3613 3427 3627
rect 3433 3613 3447 3627
rect 3393 3553 3407 3567
rect 3413 3533 3427 3547
rect 3433 3533 3447 3547
rect 3393 3493 3407 3507
rect 3433 3493 3447 3507
rect 3293 3473 3307 3487
rect 3293 3393 3307 3407
rect 3273 3293 3287 3307
rect 3213 3273 3227 3287
rect 3133 3253 3147 3267
rect 3013 3233 3027 3247
rect 3033 3213 3047 3227
rect 3053 3233 3067 3247
rect 3093 3233 3107 3247
rect 3033 3193 3047 3207
rect 3113 3213 3127 3227
rect 3133 3213 3147 3227
rect 3153 3233 3167 3247
rect 3233 3213 3247 3227
rect 3093 3193 3107 3207
rect 3173 3193 3187 3207
rect 3073 3173 3087 3187
rect 3053 3053 3067 3067
rect 3033 3033 3047 3047
rect 3113 3073 3127 3087
rect 3153 3073 3167 3087
rect 3093 3053 3107 3067
rect 3073 3033 3087 3047
rect 2993 2993 3007 3007
rect 3033 2993 3047 3007
rect 2973 2973 2987 2987
rect 2993 2853 3007 2867
rect 2953 2833 2967 2847
rect 2913 2773 2927 2787
rect 2873 2713 2887 2727
rect 2713 2693 2727 2707
rect 2793 2693 2807 2707
rect 2633 2673 2647 2687
rect 2693 2593 2707 2607
rect 2573 2513 2587 2527
rect 2553 2493 2567 2507
rect 2573 2493 2587 2507
rect 2513 2333 2527 2347
rect 2353 2293 2367 2307
rect 2393 2293 2407 2307
rect 2293 2253 2307 2267
rect 2313 2253 2327 2267
rect 2373 2273 2387 2287
rect 2273 2233 2287 2247
rect 2353 2233 2367 2247
rect 2373 2233 2387 2247
rect 2253 2213 2267 2227
rect 2233 2153 2247 2167
rect 2213 2113 2227 2127
rect 2073 1933 2087 1947
rect 2093 1933 2107 1947
rect 2153 1933 2167 1947
rect 2073 1813 2087 1827
rect 2033 1633 2047 1647
rect 2013 1613 2027 1627
rect 2233 1973 2247 1987
rect 2193 1853 2207 1867
rect 2153 1833 2167 1847
rect 2133 1773 2147 1787
rect 2193 1813 2207 1827
rect 2293 2133 2307 2147
rect 2273 2093 2287 2107
rect 2273 1833 2287 1847
rect 2173 1793 2187 1807
rect 2153 1633 2167 1647
rect 2193 1773 2207 1787
rect 2253 1793 2267 1807
rect 2273 1793 2287 1807
rect 2153 1613 2167 1627
rect 2173 1613 2187 1627
rect 2213 1753 2227 1767
rect 2013 1593 2027 1607
rect 2093 1593 2107 1607
rect 1973 1553 1987 1567
rect 1993 1553 2007 1567
rect 2053 1573 2067 1587
rect 2033 1553 2047 1567
rect 2113 1573 2127 1587
rect 2193 1593 2207 1607
rect 2333 2053 2347 2067
rect 2513 2293 2527 2307
rect 2413 2253 2427 2267
rect 2433 2273 2447 2287
rect 2473 2273 2487 2287
rect 2533 2273 2547 2287
rect 2553 2293 2567 2307
rect 2673 2553 2687 2567
rect 2693 2533 2707 2547
rect 2833 2573 2847 2587
rect 2853 2573 2867 2587
rect 2893 2573 2907 2587
rect 2733 2553 2747 2567
rect 2793 2553 2807 2567
rect 2773 2533 2787 2547
rect 2793 2513 2807 2527
rect 2853 2513 2867 2527
rect 2653 2493 2667 2507
rect 2713 2493 2727 2507
rect 2813 2493 2827 2507
rect 2873 2493 2887 2507
rect 2633 2353 2647 2367
rect 2613 2313 2627 2327
rect 2673 2333 2687 2347
rect 2613 2293 2627 2307
rect 2573 2253 2587 2267
rect 2453 2193 2467 2207
rect 2393 2093 2407 2107
rect 2413 2053 2427 2067
rect 2533 2233 2547 2247
rect 2613 2233 2627 2247
rect 2533 2153 2547 2167
rect 2593 2153 2607 2167
rect 2373 1973 2387 1987
rect 2513 1953 2527 1967
rect 2393 1933 2407 1947
rect 2393 1853 2407 1867
rect 2353 1833 2367 1847
rect 2333 1813 2347 1827
rect 2333 1793 2347 1807
rect 2373 1793 2387 1807
rect 2293 1713 2307 1727
rect 2233 1573 2247 1587
rect 2093 1553 2107 1567
rect 2173 1553 2187 1567
rect 2353 1733 2367 1747
rect 2353 1633 2367 1647
rect 2113 1533 2127 1547
rect 2333 1553 2347 1567
rect 2053 1373 2067 1387
rect 2093 1373 2107 1387
rect 1993 1333 2007 1347
rect 1993 1313 2007 1327
rect 2033 1313 2047 1327
rect 1973 1273 1987 1287
rect 1933 1253 1947 1267
rect 1953 1253 1967 1267
rect 1813 1093 1827 1107
rect 1893 1093 1907 1107
rect 1873 1073 1887 1087
rect 1913 1073 1927 1087
rect 1793 1053 1807 1067
rect 1833 1053 1847 1067
rect 2013 1233 2027 1247
rect 2013 1213 2027 1227
rect 1933 1053 1947 1067
rect 1813 1033 1827 1047
rect 1793 973 1807 987
rect 1773 933 1787 947
rect 1753 853 1767 867
rect 1753 813 1767 827
rect 1773 813 1787 827
rect 1733 753 1747 767
rect 1813 953 1827 967
rect 1953 1033 1967 1047
rect 1893 1013 1907 1027
rect 1833 913 1847 927
rect 1833 873 1847 887
rect 1933 893 1947 907
rect 1933 873 1947 887
rect 2473 1833 2487 1847
rect 2413 1753 2427 1767
rect 2413 1733 2427 1747
rect 2453 1733 2467 1747
rect 2573 2093 2587 2107
rect 2553 2073 2567 2087
rect 2653 2213 2667 2227
rect 2793 2253 2807 2267
rect 2693 2193 2707 2207
rect 2673 2153 2687 2167
rect 2653 2133 2667 2147
rect 2673 2073 2687 2087
rect 2673 2033 2687 2047
rect 2713 2053 2727 2067
rect 2733 2033 2747 2047
rect 2753 2033 2767 2047
rect 2773 2053 2787 2067
rect 2793 2033 2807 2047
rect 2613 1993 2627 2007
rect 2693 1993 2707 2007
rect 2653 1973 2667 1987
rect 2493 1773 2507 1787
rect 2533 1773 2547 1787
rect 2493 1753 2507 1767
rect 2473 1673 2487 1687
rect 2433 1633 2447 1647
rect 2433 1613 2447 1627
rect 2373 1533 2387 1547
rect 2153 1313 2167 1327
rect 2173 1313 2187 1327
rect 2193 1333 2207 1347
rect 2153 1293 2167 1307
rect 2073 1273 2087 1287
rect 2133 1273 2147 1287
rect 2093 1253 2107 1267
rect 2053 1133 2067 1147
rect 2133 1233 2147 1247
rect 2113 1093 2127 1107
rect 2133 1113 2147 1127
rect 2273 1333 2287 1347
rect 2353 1333 2367 1347
rect 2253 1293 2267 1307
rect 2333 1293 2347 1307
rect 2213 1233 2227 1247
rect 2213 1133 2227 1147
rect 2153 1093 2167 1107
rect 2073 1073 2087 1087
rect 2173 1073 2187 1087
rect 2193 1093 2207 1107
rect 2353 1133 2367 1147
rect 2033 1053 2047 1067
rect 2273 1073 2287 1087
rect 2373 1093 2387 1107
rect 2393 1113 2407 1127
rect 2253 1053 2267 1067
rect 2313 1053 2327 1067
rect 2013 1013 2027 1027
rect 1993 873 2007 887
rect 1873 853 1887 867
rect 1813 813 1827 827
rect 1793 793 1807 807
rect 1853 773 1867 787
rect 1833 753 1847 767
rect 1753 733 1767 747
rect 1593 673 1607 687
rect 1593 653 1607 667
rect 1653 653 1667 667
rect 1593 613 1607 627
rect 1733 673 1747 687
rect 1713 653 1727 667
rect 1573 593 1587 607
rect 1393 453 1407 467
rect 1353 413 1367 427
rect 1373 413 1387 427
rect 1253 373 1267 387
rect 1273 373 1287 387
rect 1333 373 1347 387
rect 1133 353 1147 367
rect 993 313 1007 327
rect 1053 313 1067 327
rect 953 193 967 207
rect 1033 293 1047 307
rect 1013 213 1027 227
rect 1153 333 1167 347
rect 1233 333 1247 347
rect 1253 333 1267 347
rect 1313 353 1327 367
rect 1113 313 1127 327
rect 1173 313 1187 327
rect 1133 293 1147 307
rect 1093 213 1107 227
rect 1113 213 1127 227
rect 1033 193 1047 207
rect 1073 193 1087 207
rect 973 173 987 187
rect 993 173 1007 187
rect 913 153 927 167
rect 933 133 947 147
rect 1253 293 1267 307
rect 1193 273 1207 287
rect 1273 233 1287 247
rect 1213 193 1227 207
rect 973 133 987 147
rect 1053 133 1067 147
rect 1093 153 1107 167
rect 1113 133 1127 147
rect 1193 133 1207 147
rect 873 113 887 127
rect 993 113 1007 127
rect 973 73 987 87
rect 1453 393 1467 407
rect 1353 353 1367 367
rect 1393 353 1407 367
rect 1333 273 1347 287
rect 1413 333 1427 347
rect 1473 333 1487 347
rect 1413 313 1427 327
rect 1373 253 1387 267
rect 1393 253 1407 267
rect 1453 313 1467 327
rect 1473 313 1487 327
rect 1433 273 1447 287
rect 1373 233 1387 247
rect 1413 233 1427 247
rect 1293 193 1307 207
rect 1313 173 1327 187
rect 1233 133 1247 147
rect 1253 113 1267 127
rect 1293 113 1307 127
rect 1213 53 1227 67
rect 853 33 867 47
rect 1333 153 1347 167
rect 1433 173 1447 187
rect 1493 293 1507 307
rect 1473 253 1487 267
rect 1533 513 1547 527
rect 1553 513 1567 527
rect 1773 653 1787 667
rect 1813 653 1827 667
rect 1753 613 1767 627
rect 1673 573 1687 587
rect 1653 533 1667 547
rect 1593 513 1607 527
rect 1633 513 1647 527
rect 1593 433 1607 447
rect 1553 373 1567 387
rect 1573 373 1587 387
rect 1533 353 1547 367
rect 1533 273 1547 287
rect 1633 393 1647 407
rect 1653 393 1667 407
rect 1713 593 1727 607
rect 1753 593 1767 607
rect 1773 573 1787 587
rect 1693 513 1707 527
rect 1733 493 1747 507
rect 1713 473 1727 487
rect 1693 413 1707 427
rect 1713 413 1727 427
rect 1673 373 1687 387
rect 1973 853 1987 867
rect 1913 793 1927 807
rect 1953 793 1967 807
rect 1933 773 1947 787
rect 1873 673 1887 687
rect 1833 593 1847 607
rect 1813 533 1827 547
rect 1853 573 1867 587
rect 1893 573 1907 587
rect 1833 513 1847 527
rect 1833 493 1847 507
rect 1773 473 1787 487
rect 1793 473 1807 487
rect 1813 393 1827 407
rect 1633 353 1647 367
rect 1673 353 1687 367
rect 1593 273 1607 287
rect 1573 253 1587 267
rect 1713 353 1727 367
rect 1753 353 1767 367
rect 1733 333 1747 347
rect 1673 313 1687 327
rect 1693 313 1707 327
rect 1653 253 1667 267
rect 1633 233 1647 247
rect 1693 293 1707 307
rect 1753 293 1767 307
rect 1533 193 1547 207
rect 1613 193 1627 207
rect 1493 173 1507 187
rect 1513 173 1527 187
rect 1433 153 1447 167
rect 1353 113 1367 127
rect 1433 133 1447 147
rect 1473 133 1487 147
rect 1553 153 1567 167
rect 1533 133 1547 147
rect 1513 113 1527 127
rect 1573 133 1587 147
rect 1613 133 1627 147
rect 1693 233 1707 247
rect 1673 173 1687 187
rect 1693 173 1707 187
rect 1733 173 1747 187
rect 1873 453 1887 467
rect 1913 453 1927 467
rect 1853 433 1867 447
rect 1913 433 1927 447
rect 1893 413 1907 427
rect 1913 393 1927 407
rect 2153 933 2167 947
rect 2053 833 2067 847
rect 2013 793 2027 807
rect 1993 773 2007 787
rect 1993 753 2007 767
rect 1973 733 1987 747
rect 1953 713 1967 727
rect 2053 773 2067 787
rect 2033 713 2047 727
rect 2013 653 2027 667
rect 2053 693 2067 707
rect 2133 833 2147 847
rect 2093 693 2107 707
rect 1993 613 2007 627
rect 2133 733 2147 747
rect 2113 653 2127 667
rect 2113 633 2127 647
rect 2093 613 2107 627
rect 1973 593 1987 607
rect 2013 533 2027 547
rect 2033 533 2047 547
rect 1993 473 2007 487
rect 1953 393 1967 407
rect 2113 593 2127 607
rect 2093 553 2107 567
rect 2053 513 2067 527
rect 2033 413 2047 427
rect 2173 813 2187 827
rect 2193 833 2207 847
rect 2213 813 2227 827
rect 2513 1733 2527 1747
rect 2593 1793 2607 1807
rect 2633 1793 2647 1807
rect 2673 1953 2687 1967
rect 2753 1993 2767 2007
rect 2733 1833 2747 1847
rect 2573 1753 2587 1767
rect 2553 1673 2567 1687
rect 2553 1653 2567 1667
rect 2733 1813 2747 1827
rect 2693 1773 2707 1787
rect 2853 2273 2867 2287
rect 2913 2553 2927 2567
rect 2973 2733 2987 2747
rect 3013 2713 3027 2727
rect 3053 2973 3067 2987
rect 3033 2673 3047 2687
rect 2993 2633 3007 2647
rect 3033 2573 3047 2587
rect 2913 2513 2927 2527
rect 2933 2533 2947 2547
rect 2953 2493 2967 2507
rect 2913 2413 2927 2427
rect 2973 2413 2987 2427
rect 2893 2173 2907 2187
rect 3533 3733 3547 3747
rect 3573 3733 3587 3747
rect 3553 3693 3567 3707
rect 3713 3713 3727 3727
rect 3733 3693 3747 3707
rect 3693 3673 3707 3687
rect 3633 3633 3647 3647
rect 3493 3593 3507 3607
rect 3593 3593 3607 3607
rect 3473 3553 3487 3567
rect 3473 3533 3487 3547
rect 3533 3553 3547 3567
rect 3573 3553 3587 3567
rect 3513 3533 3527 3547
rect 3553 3493 3567 3507
rect 3613 3513 3627 3527
rect 3493 3473 3507 3487
rect 3553 3473 3567 3487
rect 3473 3333 3487 3347
rect 3473 3313 3487 3327
rect 3433 3253 3447 3267
rect 3293 3233 3307 3247
rect 3273 3193 3287 3207
rect 3253 3113 3267 3127
rect 3213 3053 3227 3067
rect 3153 3013 3167 3027
rect 3173 3013 3187 3027
rect 3193 3033 3207 3047
rect 3133 2993 3147 3007
rect 3093 2933 3107 2947
rect 3093 2873 3107 2887
rect 3093 2793 3107 2807
rect 3113 2693 3127 2707
rect 3253 2973 3267 2987
rect 3253 2713 3267 2727
rect 3213 2693 3227 2707
rect 3313 3213 3327 3227
rect 3353 3233 3367 3247
rect 3373 3213 3387 3227
rect 3453 3213 3467 3227
rect 3333 3153 3347 3167
rect 3393 3193 3407 3207
rect 3393 3093 3407 3107
rect 3293 2993 3307 3007
rect 3213 2673 3227 2687
rect 3153 2653 3167 2667
rect 3073 2553 3087 2567
rect 3093 2533 3107 2547
rect 3133 2533 3147 2547
rect 3093 2353 3107 2367
rect 2993 2293 3007 2307
rect 2933 2253 2947 2267
rect 2933 2233 2947 2247
rect 2913 2153 2927 2167
rect 2913 2073 2927 2087
rect 2973 2253 2987 2267
rect 2953 2193 2967 2207
rect 2973 2173 2987 2187
rect 3013 2173 3027 2187
rect 2913 2033 2927 2047
rect 2813 1933 2827 1947
rect 2773 1773 2787 1787
rect 2853 1793 2867 1807
rect 2893 1793 2907 1807
rect 2933 1853 2947 1867
rect 2953 1793 2967 1807
rect 2873 1773 2887 1787
rect 2913 1773 2927 1787
rect 2793 1753 2807 1767
rect 2813 1753 2827 1767
rect 2833 1753 2847 1767
rect 2773 1673 2787 1687
rect 2613 1633 2627 1647
rect 2673 1633 2687 1647
rect 2713 1633 2727 1647
rect 2753 1633 2767 1647
rect 2593 1613 2607 1627
rect 2533 1593 2547 1607
rect 2533 1573 2547 1587
rect 2573 1573 2587 1587
rect 2733 1613 2747 1627
rect 2833 1673 2847 1687
rect 2933 1633 2947 1647
rect 2633 1593 2647 1607
rect 2693 1593 2707 1607
rect 2833 1613 2847 1627
rect 2933 1613 2947 1627
rect 2753 1593 2767 1607
rect 2793 1573 2807 1587
rect 2833 1573 2847 1587
rect 2853 1593 2867 1607
rect 2893 1593 2907 1607
rect 2913 1593 2927 1607
rect 2873 1573 2887 1587
rect 2553 1553 2567 1567
rect 2613 1553 2627 1567
rect 2653 1553 2667 1567
rect 2773 1553 2787 1567
rect 2493 1493 2507 1507
rect 2433 1333 2447 1347
rect 2473 1333 2487 1347
rect 2513 1313 2527 1327
rect 2793 1533 2807 1547
rect 2653 1353 2667 1367
rect 2593 1333 2607 1347
rect 2713 1333 2727 1347
rect 2813 1333 2827 1347
rect 2593 1293 2607 1307
rect 2633 1293 2647 1307
rect 2673 1293 2687 1307
rect 2753 1293 2767 1307
rect 2773 1313 2787 1327
rect 2813 1313 2827 1327
rect 2833 1293 2847 1307
rect 2453 1273 2467 1287
rect 2493 1273 2507 1287
rect 2793 1233 2807 1247
rect 2693 1193 2707 1207
rect 2633 1173 2647 1187
rect 2453 1093 2467 1107
rect 2613 1133 2627 1147
rect 2673 1153 2687 1167
rect 2853 1173 2867 1187
rect 2693 1133 2707 1147
rect 2593 1113 2607 1127
rect 2513 1073 2527 1087
rect 2533 1093 2547 1107
rect 2613 1093 2627 1107
rect 2653 1093 2667 1107
rect 2733 1113 2747 1127
rect 2793 1113 2807 1127
rect 2553 1073 2567 1087
rect 2653 1073 2667 1087
rect 2513 973 2527 987
rect 2493 953 2507 967
rect 2413 873 2427 887
rect 2353 853 2367 867
rect 2273 813 2287 827
rect 2313 833 2327 847
rect 2393 833 2407 847
rect 2433 833 2447 847
rect 2173 793 2187 807
rect 2233 793 2247 807
rect 2293 793 2307 807
rect 2253 773 2267 787
rect 2193 753 2207 767
rect 2153 593 2167 607
rect 2173 613 2187 627
rect 2233 673 2247 687
rect 2273 733 2287 747
rect 2433 753 2447 767
rect 2373 693 2387 707
rect 2333 673 2347 687
rect 2373 673 2387 687
rect 2313 653 2327 667
rect 2333 653 2347 667
rect 2413 653 2427 667
rect 2213 633 2227 647
rect 2253 633 2267 647
rect 2193 593 2207 607
rect 2173 573 2187 587
rect 2173 533 2187 547
rect 2133 513 2147 527
rect 2133 473 2147 487
rect 2173 473 2187 487
rect 2113 413 2127 427
rect 2193 453 2207 467
rect 1933 373 1947 387
rect 1873 353 1887 367
rect 1813 333 1827 347
rect 1833 333 1847 347
rect 1793 273 1807 287
rect 1773 253 1787 267
rect 1773 193 1787 207
rect 1753 153 1767 167
rect 1673 133 1687 147
rect 1693 133 1707 147
rect 1733 133 1747 147
rect 1593 113 1607 127
rect 1633 113 1647 127
rect 1393 93 1407 107
rect 1473 73 1487 87
rect 1313 13 1327 27
rect 1713 113 1727 127
rect 1753 113 1767 127
rect 1913 333 1927 347
rect 1853 313 1867 327
rect 1873 253 1887 267
rect 1913 153 1927 167
rect 1813 113 1827 127
rect 1893 113 1907 127
rect 1913 113 1927 127
rect 1693 93 1707 107
rect 1793 93 1807 107
rect 1833 73 1847 87
rect 1513 53 1527 67
rect 1753 53 1767 67
rect 1873 33 1887 47
rect 1913 73 1927 87
rect 1993 373 2007 387
rect 2013 353 2027 367
rect 2053 353 2067 367
rect 2073 373 2087 387
rect 2093 373 2107 387
rect 1953 293 1967 307
rect 2053 333 2067 347
rect 2133 353 2147 367
rect 2013 313 2027 327
rect 1993 293 2007 307
rect 2033 293 2047 307
rect 1973 253 1987 267
rect 1953 173 1967 187
rect 1973 153 1987 167
rect 1933 33 1947 47
rect 2013 213 2027 227
rect 2073 233 2087 247
rect 2093 193 2107 207
rect 2053 173 2067 187
rect 2073 173 2087 187
rect 2013 153 2027 167
rect 1993 93 2007 107
rect 2053 73 2067 87
rect 2133 293 2147 307
rect 2213 373 2227 387
rect 2293 613 2307 627
rect 2353 613 2367 627
rect 2393 633 2407 647
rect 2273 593 2287 607
rect 2293 593 2307 607
rect 2493 853 2507 867
rect 2453 693 2467 707
rect 2473 673 2487 687
rect 2553 953 2567 967
rect 2953 1593 2967 1607
rect 2893 1553 2907 1567
rect 2913 1533 2927 1547
rect 2873 1153 2887 1167
rect 2893 1153 2907 1167
rect 2993 2113 3007 2127
rect 3193 2553 3207 2567
rect 3153 2293 3167 2307
rect 3053 2253 3067 2267
rect 3073 2253 3087 2267
rect 3173 2253 3187 2267
rect 3193 2253 3207 2267
rect 3113 2193 3127 2207
rect 3033 2113 3047 2127
rect 3053 2093 3067 2107
rect 3233 2593 3247 2607
rect 3373 3073 3387 3087
rect 3533 3333 3547 3347
rect 3533 3253 3547 3267
rect 3473 3193 3487 3207
rect 3353 3033 3367 3047
rect 3433 3033 3447 3047
rect 3393 2993 3407 3007
rect 3493 3073 3507 3087
rect 3493 3013 3507 3027
rect 3373 2953 3387 2967
rect 3293 2613 3307 2627
rect 3333 2573 3347 2587
rect 3353 2573 3367 2587
rect 3433 2933 3447 2947
rect 3593 3313 3607 3327
rect 3653 3573 3667 3587
rect 3673 3553 3687 3567
rect 3653 3533 3667 3547
rect 3813 4193 3827 4207
rect 3833 4193 3847 4207
rect 3973 4513 3987 4527
rect 3953 4373 3967 4387
rect 3933 4213 3947 4227
rect 3873 4173 3887 4187
rect 3913 4173 3927 4187
rect 3913 4133 3927 4147
rect 3873 4073 3887 4087
rect 3853 4033 3867 4047
rect 3933 4033 3947 4047
rect 3813 3993 3827 4007
rect 3913 4013 3927 4027
rect 3833 3973 3847 3987
rect 3853 3973 3867 3987
rect 3893 3993 3907 4007
rect 4053 4573 4067 4587
rect 4033 4553 4047 4567
rect 4113 4573 4127 4587
rect 4133 4573 4147 4587
rect 4153 4553 4167 4567
rect 4233 4573 4247 4587
rect 4193 4533 4207 4547
rect 4133 4493 4147 4507
rect 4153 4493 4167 4507
rect 4113 4473 4127 4487
rect 4093 4433 4107 4447
rect 4173 4433 4187 4447
rect 4053 4413 4067 4427
rect 4033 4393 4047 4407
rect 4233 4453 4247 4467
rect 4193 4393 4207 4407
rect 4033 4293 4047 4307
rect 4093 4293 4107 4307
rect 4133 4293 4147 4307
rect 4013 4153 4027 4167
rect 4193 4233 4207 4247
rect 4213 4233 4227 4247
rect 4133 4213 4147 4227
rect 4053 4173 4067 4187
rect 4173 4193 4187 4207
rect 4073 4153 4087 4167
rect 4033 4093 4047 4107
rect 4193 4153 4207 4167
rect 4313 4573 4327 4587
rect 4353 4573 4367 4587
rect 4333 4493 4347 4507
rect 4273 4473 4287 4487
rect 4293 4453 4307 4467
rect 4313 4473 4327 4487
rect 4293 4433 4307 4447
rect 4273 4173 4287 4187
rect 4213 4093 4227 4107
rect 4233 4093 4247 4107
rect 4033 4053 4047 4067
rect 4073 4053 4087 4067
rect 4093 4053 4107 4067
rect 4133 4053 4147 4067
rect 4193 4053 4207 4067
rect 3853 3933 3867 3947
rect 3813 3913 3827 3927
rect 3873 3913 3887 3927
rect 3773 3673 3787 3687
rect 3793 3673 3807 3687
rect 3813 3653 3827 3667
rect 3893 3713 3907 3727
rect 3873 3693 3887 3707
rect 3813 3593 3827 3607
rect 3753 3533 3767 3547
rect 3713 3493 3727 3507
rect 3753 3493 3767 3507
rect 3793 3493 3807 3507
rect 3853 3513 3867 3527
rect 3693 3473 3707 3487
rect 3773 3453 3787 3467
rect 3833 3453 3847 3467
rect 3833 3433 3847 3447
rect 3573 3293 3587 3307
rect 3593 3293 3607 3307
rect 3633 3293 3647 3307
rect 3593 3233 3607 3247
rect 3613 3253 3627 3267
rect 3773 3313 3787 3327
rect 3693 3253 3707 3267
rect 3573 3133 3587 3147
rect 3633 3133 3647 3147
rect 3533 3013 3547 3027
rect 3413 2713 3427 2727
rect 3433 2713 3447 2727
rect 3493 2733 3507 2747
rect 3453 2673 3467 2687
rect 3493 2693 3507 2707
rect 3453 2633 3467 2647
rect 3473 2633 3487 2647
rect 3473 2593 3487 2607
rect 3293 2533 3307 2547
rect 3393 2533 3407 2547
rect 3473 2553 3487 2567
rect 3313 2513 3327 2527
rect 3273 2493 3287 2507
rect 3253 2453 3267 2467
rect 3293 2313 3307 2327
rect 3233 2253 3247 2267
rect 3253 2253 3267 2267
rect 3213 2213 3227 2227
rect 3133 2173 3147 2187
rect 3173 2173 3187 2187
rect 3093 2073 3107 2087
rect 3193 2113 3207 2127
rect 3213 2093 3227 2107
rect 3133 2053 3147 2067
rect 3153 2053 3167 2067
rect 3173 2073 3187 2087
rect 3113 2033 3127 2047
rect 3133 1993 3147 2007
rect 3153 1853 3167 1867
rect 3053 1813 3067 1827
rect 3053 1773 3067 1787
rect 3073 1773 3087 1787
rect 3093 1773 3107 1787
rect 3033 1753 3047 1767
rect 3133 1813 3147 1827
rect 3133 1693 3147 1707
rect 3133 1633 3147 1647
rect 3213 1633 3227 1647
rect 2993 1613 3007 1627
rect 2993 1573 3007 1587
rect 3333 2233 3347 2247
rect 3393 2513 3407 2527
rect 3433 2513 3447 2527
rect 3373 2253 3387 2267
rect 3353 2213 3367 2227
rect 3293 2193 3307 2207
rect 3253 2153 3267 2167
rect 3273 2133 3287 2147
rect 3253 2053 3267 2067
rect 3293 2053 3307 2067
rect 3313 2073 3327 2087
rect 3333 2053 3347 2067
rect 3273 1933 3287 1947
rect 3253 1693 3267 1707
rect 3053 1573 3067 1587
rect 3093 1593 3107 1607
rect 3113 1573 3127 1587
rect 3173 1593 3187 1607
rect 3233 1593 3247 1607
rect 3153 1573 3167 1587
rect 3213 1573 3227 1587
rect 3233 1553 3247 1567
rect 3173 1533 3187 1547
rect 3193 1533 3207 1547
rect 2973 1353 2987 1367
rect 2993 1313 3007 1327
rect 2973 1273 2987 1287
rect 2933 1253 2947 1267
rect 2973 1153 2987 1167
rect 2993 1133 3007 1147
rect 2973 1113 2987 1127
rect 3253 1373 3267 1387
rect 3173 1353 3187 1367
rect 3253 1353 3267 1367
rect 3093 1333 3107 1347
rect 3053 1293 3067 1307
rect 3073 1293 3087 1307
rect 3013 1113 3027 1127
rect 3033 1093 3047 1107
rect 3113 1293 3127 1307
rect 3213 1333 3227 1347
rect 3193 1253 3207 1267
rect 3233 1253 3247 1267
rect 3373 2033 3387 2047
rect 3453 2073 3467 2087
rect 3433 2013 3447 2027
rect 3293 1833 3307 1847
rect 3333 1833 3347 1847
rect 3453 1833 3467 1847
rect 3333 1793 3347 1807
rect 3373 1793 3387 1807
rect 3413 1813 3427 1827
rect 3433 1793 3447 1807
rect 3373 1773 3387 1787
rect 3353 1733 3367 1747
rect 3333 1653 3347 1667
rect 3313 1633 3327 1647
rect 3353 1613 3367 1627
rect 3333 1593 3347 1607
rect 3333 1553 3347 1567
rect 3333 1533 3347 1547
rect 3293 1513 3307 1527
rect 3293 1373 3307 1387
rect 3273 1193 3287 1207
rect 3133 1153 3147 1167
rect 3173 1133 3187 1147
rect 3213 1133 3227 1147
rect 2913 1053 2927 1067
rect 3113 1093 3127 1107
rect 3253 1113 3267 1127
rect 2993 1053 3007 1067
rect 2553 853 2567 867
rect 2753 853 2767 867
rect 2573 833 2587 847
rect 2593 833 2607 847
rect 2633 833 2647 847
rect 2573 793 2587 807
rect 2613 813 2627 827
rect 2673 833 2687 847
rect 2773 833 2787 847
rect 2793 853 2807 867
rect 2893 853 2907 867
rect 2933 853 2947 867
rect 2693 813 2707 827
rect 2833 813 2847 827
rect 2853 833 2867 847
rect 2913 813 2927 827
rect 2653 793 2667 807
rect 2573 733 2587 747
rect 2533 713 2547 727
rect 2453 653 2467 667
rect 2513 653 2527 667
rect 2473 633 2487 647
rect 2453 613 2467 627
rect 2473 613 2487 627
rect 2453 593 2467 607
rect 2513 613 2527 627
rect 2493 593 2507 607
rect 2413 493 2427 507
rect 2293 473 2307 487
rect 2273 433 2287 447
rect 2413 413 2427 427
rect 2333 393 2347 407
rect 2193 353 2207 367
rect 2233 353 2247 367
rect 2333 373 2347 387
rect 2273 333 2287 347
rect 2313 333 2327 347
rect 2353 333 2367 347
rect 2213 313 2227 327
rect 2193 273 2207 287
rect 2133 213 2147 227
rect 2173 213 2187 227
rect 2193 213 2207 227
rect 2153 193 2167 207
rect 2173 193 2187 207
rect 2113 53 2127 67
rect 2213 153 2227 167
rect 2373 313 2387 327
rect 2253 293 2267 307
rect 2393 293 2407 307
rect 2253 273 2267 287
rect 2393 253 2407 267
rect 2253 193 2267 207
rect 2353 193 2367 207
rect 2353 173 2367 187
rect 2433 353 2447 367
rect 2433 333 2447 347
rect 2413 193 2427 207
rect 2493 373 2507 387
rect 2473 333 2487 347
rect 2453 213 2467 227
rect 2553 593 2567 607
rect 2673 653 2687 667
rect 2693 633 2707 647
rect 2773 633 2787 647
rect 2673 613 2687 627
rect 2653 593 2667 607
rect 2733 613 2747 627
rect 2713 593 2727 607
rect 2673 533 2687 547
rect 2733 533 2747 547
rect 2553 413 2567 427
rect 2633 413 2647 427
rect 2533 373 2547 387
rect 2573 393 2587 407
rect 2693 393 2707 407
rect 2573 353 2587 367
rect 2633 353 2647 367
rect 2533 293 2547 307
rect 2553 193 2567 207
rect 2593 173 2607 187
rect 2173 133 2187 147
rect 2193 133 2207 147
rect 2313 153 2327 167
rect 2333 133 2347 147
rect 2413 133 2427 147
rect 2753 393 2767 407
rect 2733 373 2747 387
rect 2913 713 2927 727
rect 2953 833 2967 847
rect 2973 793 2987 807
rect 3073 833 3087 847
rect 3053 813 3067 827
rect 3013 793 3027 807
rect 2993 753 3007 767
rect 2953 713 2967 727
rect 2933 633 2947 647
rect 2873 413 2887 427
rect 2853 373 2867 387
rect 2673 353 2687 367
rect 2773 353 2787 367
rect 2753 333 2767 347
rect 2793 333 2807 347
rect 2653 313 2667 327
rect 2713 313 2727 327
rect 2833 333 2847 347
rect 2893 373 2907 387
rect 2913 353 2927 367
rect 2933 373 2947 387
rect 2873 333 2887 347
rect 2813 313 2827 327
rect 2853 313 2867 327
rect 2653 253 2667 267
rect 2693 253 2707 267
rect 2253 113 2267 127
rect 2233 93 2247 107
rect 2573 133 2587 147
rect 2593 153 2607 167
rect 3093 793 3107 807
rect 3153 793 3167 807
rect 3233 833 3247 847
rect 3253 813 3267 827
rect 3073 773 3087 787
rect 3113 773 3127 787
rect 3133 773 3147 787
rect 3193 773 3207 787
rect 3073 753 3087 767
rect 3033 653 3047 667
rect 3193 653 3207 667
rect 3213 653 3227 667
rect 3233 653 3247 667
rect 3273 653 3287 667
rect 3173 633 3187 647
rect 3093 613 3107 627
rect 3153 613 3167 627
rect 3053 593 3067 607
rect 3013 373 3027 387
rect 2973 293 2987 307
rect 2713 133 2727 147
rect 2533 113 2547 127
rect 2613 113 2627 127
rect 2473 93 2487 107
rect 2953 233 2967 247
rect 2773 193 2787 207
rect 2853 173 2867 187
rect 2773 153 2787 167
rect 2753 133 2767 147
rect 2793 133 2807 147
rect 2873 133 2887 147
rect 2293 73 2307 87
rect 2733 73 2747 87
rect 2813 73 2827 87
rect 3013 233 3027 247
rect 3453 1753 3467 1767
rect 3393 1613 3407 1627
rect 3373 1573 3387 1587
rect 3433 1593 3447 1607
rect 3413 1553 3427 1567
rect 3353 1513 3367 1527
rect 3353 1233 3367 1247
rect 3533 2773 3547 2787
rect 3553 2773 3567 2787
rect 3533 2653 3547 2667
rect 3533 2613 3547 2627
rect 3513 2513 3527 2527
rect 3633 3093 3647 3107
rect 3753 3213 3767 3227
rect 3913 3573 3927 3587
rect 4013 4013 4027 4027
rect 3993 3993 4007 4007
rect 4053 3993 4067 4007
rect 3973 3953 3987 3967
rect 4093 4033 4107 4047
rect 4113 3993 4127 4007
rect 4153 4013 4167 4027
rect 4173 3973 4187 3987
rect 4193 3993 4207 4007
rect 4213 3973 4227 3987
rect 4053 3833 4067 3847
rect 3913 3533 3927 3547
rect 3953 3533 3967 3547
rect 3953 3513 3967 3527
rect 3893 3453 3907 3467
rect 3933 3453 3947 3467
rect 3873 3393 3887 3407
rect 4233 3853 4247 3867
rect 4393 4393 4407 4407
rect 4353 4213 4367 4227
rect 4313 4193 4327 4207
rect 4373 4173 4387 4187
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4333 4153 4347 4167
rect 4453 4153 4467 4167
rect 4513 4473 4527 4487
rect 4553 4233 4567 4247
rect 4513 4173 4527 4187
rect 4493 4133 4507 4147
rect 4513 4133 4527 4147
rect 4373 4113 4387 4127
rect 4413 4113 4427 4127
rect 4293 4093 4307 4107
rect 4273 4073 4287 4087
rect 4333 4073 4347 4087
rect 4273 3993 4287 4007
rect 4293 3993 4307 4007
rect 4313 3973 4327 3987
rect 4413 3973 4427 3987
rect 4293 3853 4307 3867
rect 4253 3733 4267 3747
rect 4073 3673 4087 3687
rect 4053 3573 4067 3587
rect 4033 3553 4047 3567
rect 4033 3533 4047 3547
rect 4013 3453 4027 3467
rect 3893 3273 3907 3287
rect 3913 3273 3927 3287
rect 3953 3273 3967 3287
rect 3973 3273 3987 3287
rect 4013 3273 4027 3287
rect 3873 3253 3887 3267
rect 3813 3153 3827 3167
rect 3833 3153 3847 3167
rect 3713 3093 3727 3107
rect 3673 3053 3687 3067
rect 3633 3033 3647 3047
rect 3673 3033 3687 3047
rect 3613 3013 3627 3027
rect 3653 2993 3667 3007
rect 3633 2873 3647 2887
rect 3593 2773 3607 2787
rect 3593 2733 3607 2747
rect 3613 2633 3627 2647
rect 3593 2553 3607 2567
rect 3553 2493 3567 2507
rect 3573 2493 3587 2507
rect 3533 2353 3547 2367
rect 3573 2353 3587 2367
rect 3553 2293 3567 2307
rect 3493 2273 3507 2287
rect 3513 2253 3527 2267
rect 3713 3073 3727 3087
rect 3773 3073 3787 3087
rect 3713 3033 3727 3047
rect 3753 3033 3767 3047
rect 3793 3033 3807 3047
rect 3773 3013 3787 3027
rect 3813 3013 3827 3027
rect 3713 2993 3727 3007
rect 3713 2973 3727 2987
rect 3673 2853 3687 2867
rect 3653 2773 3667 2787
rect 3653 2733 3667 2747
rect 3673 2593 3687 2607
rect 3693 2553 3707 2567
rect 3673 2353 3687 2367
rect 3693 2353 3707 2367
rect 3633 2313 3647 2327
rect 3653 2313 3667 2327
rect 3493 2233 3507 2247
rect 3513 2213 3527 2227
rect 3493 2013 3507 2027
rect 3613 2273 3627 2287
rect 3593 2253 3607 2267
rect 3653 2273 3667 2287
rect 3633 2253 3647 2267
rect 3593 2233 3607 2247
rect 3673 2253 3687 2267
rect 3653 2233 3667 2247
rect 3593 2193 3607 2207
rect 3573 2173 3587 2187
rect 3533 2113 3547 2127
rect 3533 2073 3547 2087
rect 3573 2073 3587 2087
rect 3553 1853 3567 1867
rect 3513 1813 3527 1827
rect 3493 1753 3507 1767
rect 3473 1713 3487 1727
rect 3473 1593 3487 1607
rect 3473 1533 3487 1547
rect 3513 1633 3527 1647
rect 3413 1493 3427 1507
rect 3453 1493 3467 1507
rect 3393 1273 3407 1287
rect 3393 1233 3407 1247
rect 3333 1133 3347 1147
rect 3373 1193 3387 1207
rect 3373 1173 3387 1187
rect 3473 1293 3487 1307
rect 3453 1213 3467 1227
rect 3473 1153 3487 1167
rect 3413 1093 3427 1107
rect 3313 853 3327 867
rect 3333 833 3347 847
rect 3353 853 3367 867
rect 3393 853 3407 867
rect 3373 833 3387 847
rect 3413 813 3427 827
rect 3333 753 3347 767
rect 3393 753 3407 767
rect 3253 633 3267 647
rect 3293 633 3307 647
rect 3273 613 3287 627
rect 3293 613 3307 627
rect 3233 593 3247 607
rect 3353 673 3367 687
rect 3173 573 3187 587
rect 3213 573 3227 587
rect 3493 1093 3507 1107
rect 3473 813 3487 827
rect 3493 793 3507 807
rect 3493 713 3507 727
rect 3533 1613 3547 1627
rect 3673 2133 3687 2147
rect 3613 2093 3627 2107
rect 3613 2073 3627 2087
rect 3653 2073 3667 2087
rect 3633 1993 3647 2007
rect 3613 1933 3627 1947
rect 3573 1753 3587 1767
rect 3653 1853 3667 1867
rect 3573 1713 3587 1727
rect 3573 1613 3587 1627
rect 3573 1553 3587 1567
rect 3533 1313 3547 1327
rect 3553 1273 3567 1287
rect 3633 1733 3647 1747
rect 3613 1673 3627 1687
rect 3653 1633 3667 1647
rect 3813 2953 3827 2967
rect 3733 2913 3747 2927
rect 3773 2913 3787 2927
rect 3853 3113 3867 3127
rect 3913 3133 3927 3147
rect 3893 3053 3907 3067
rect 3853 3033 3867 3047
rect 3853 3013 3867 3027
rect 3893 3013 3907 3027
rect 3953 3213 3967 3227
rect 4053 3513 4067 3527
rect 4193 3713 4207 3727
rect 4233 3713 4247 3727
rect 4113 3653 4127 3667
rect 4093 3593 4107 3607
rect 4073 3433 4087 3447
rect 4073 3313 4087 3327
rect 4033 3253 4047 3267
rect 4013 3233 4027 3247
rect 3993 3213 4007 3227
rect 3973 3173 3987 3187
rect 4013 3193 4027 3207
rect 4013 3153 4027 3167
rect 3993 3133 4007 3147
rect 3993 3113 4007 3127
rect 4013 3113 4027 3127
rect 3973 3073 3987 3087
rect 4053 3153 4067 3167
rect 4093 3213 4107 3227
rect 4273 3713 4287 3727
rect 4253 3693 4267 3707
rect 4193 3673 4207 3687
rect 4173 3633 4187 3647
rect 4153 3613 4167 3627
rect 4173 3593 4187 3607
rect 4153 3553 4167 3567
rect 4153 3413 4167 3427
rect 4113 3193 4127 3207
rect 4073 3113 4087 3127
rect 4113 3093 4127 3107
rect 4013 3073 4027 3087
rect 4033 3073 4047 3087
rect 4093 3053 4107 3067
rect 3953 3033 3967 3047
rect 3993 3013 4007 3027
rect 4053 3013 4067 3027
rect 4073 3033 4087 3047
rect 4173 3233 4187 3247
rect 4213 3653 4227 3667
rect 4313 3833 4327 3847
rect 4293 3633 4307 3647
rect 4273 3613 4287 3627
rect 4313 3613 4327 3627
rect 4293 3513 4307 3527
rect 4213 3413 4227 3427
rect 4353 3593 4367 3607
rect 4373 3593 4387 3607
rect 4333 3453 4347 3467
rect 4353 3453 4367 3467
rect 4433 3693 4447 3707
rect 4553 3993 4567 4007
rect 4613 4513 4627 4527
rect 4673 4453 4687 4467
rect 4613 4433 4627 4447
rect 4593 4133 4607 4147
rect 4493 3753 4507 3767
rect 4533 3753 4547 3767
rect 4413 3613 4427 3627
rect 4413 3593 4427 3607
rect 4393 3513 4407 3527
rect 4393 3493 4407 3507
rect 4473 3513 4487 3527
rect 4453 3493 4467 3507
rect 4453 3293 4467 3307
rect 4413 3273 4427 3287
rect 4433 3273 4447 3287
rect 4493 3313 4507 3327
rect 4313 3253 4327 3267
rect 4333 3253 4347 3267
rect 4193 3213 4207 3227
rect 4233 3213 4247 3227
rect 4253 3233 4267 3247
rect 4273 3213 4287 3227
rect 4173 3173 4187 3187
rect 4213 3153 4227 3167
rect 4133 3073 4147 3087
rect 4193 3053 4207 3067
rect 4113 3013 4127 3027
rect 4173 3033 4187 3047
rect 3973 2993 3987 3007
rect 4113 2993 4127 3007
rect 4133 2993 4147 3007
rect 3833 2873 3847 2887
rect 3813 2833 3827 2847
rect 3773 2813 3787 2827
rect 3733 2693 3747 2707
rect 3793 2773 3807 2787
rect 3793 2653 3807 2667
rect 3773 2613 3787 2627
rect 3713 2313 3727 2327
rect 3713 2273 3727 2287
rect 3713 2233 3727 2247
rect 3713 1933 3727 1947
rect 3933 2813 3947 2827
rect 3853 2793 3867 2807
rect 3893 2773 3907 2787
rect 3873 2733 3887 2747
rect 3833 2713 3847 2727
rect 3773 2533 3787 2547
rect 3813 2593 3827 2607
rect 3813 2493 3827 2507
rect 3773 2393 3787 2407
rect 3813 2373 3827 2387
rect 3773 2293 3787 2307
rect 3813 2293 3827 2307
rect 3773 2253 3787 2267
rect 3753 2193 3767 2207
rect 3813 2253 3827 2267
rect 4093 2973 4107 2987
rect 4033 2813 4047 2827
rect 3973 2753 3987 2767
rect 3853 2693 3867 2707
rect 3893 2693 3907 2707
rect 3933 2693 3947 2707
rect 3913 2593 3927 2607
rect 4053 2733 4067 2747
rect 3973 2713 3987 2727
rect 4013 2713 4027 2727
rect 4053 2713 4067 2727
rect 3993 2693 4007 2707
rect 3993 2633 4007 2647
rect 4073 2693 4087 2707
rect 3973 2613 3987 2627
rect 4053 2613 4067 2627
rect 4173 2993 4187 3007
rect 4153 2953 4167 2967
rect 4133 2813 4147 2827
rect 4253 3193 4267 3207
rect 4273 3193 4287 3207
rect 4253 3153 4267 3167
rect 4253 3133 4267 3147
rect 4233 3113 4247 3127
rect 4233 3053 4247 3067
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4413 3213 4427 3227
rect 4333 3193 4347 3207
rect 4293 3133 4307 3147
rect 4293 3113 4307 3127
rect 4233 3013 4247 3027
rect 4313 3073 4327 3087
rect 4353 3173 4367 3187
rect 4393 3153 4407 3167
rect 4373 3133 4387 3147
rect 4353 3113 4367 3127
rect 4293 3033 4307 3047
rect 4293 3013 4307 3027
rect 4233 2933 4247 2947
rect 4333 3053 4347 3067
rect 4353 3033 4367 3047
rect 4353 2993 4367 3007
rect 4273 2973 4287 2987
rect 4293 2973 4307 2987
rect 4273 2913 4287 2927
rect 4273 2853 4287 2867
rect 4253 2833 4267 2847
rect 4213 2773 4227 2787
rect 4133 2753 4147 2767
rect 4113 2713 4127 2727
rect 4113 2693 4127 2707
rect 4013 2593 4027 2607
rect 4093 2593 4107 2607
rect 3953 2573 3967 2587
rect 3873 2553 3887 2567
rect 3893 2533 3907 2547
rect 3933 2533 3947 2547
rect 3953 2553 3967 2567
rect 3993 2553 4007 2567
rect 3973 2533 3987 2547
rect 3853 2473 3867 2487
rect 3933 2473 3947 2487
rect 3953 2473 3967 2487
rect 3873 2353 3887 2367
rect 4073 2573 4087 2587
rect 4033 2553 4047 2567
rect 4053 2513 4067 2527
rect 4033 2493 4047 2507
rect 4093 2493 4107 2507
rect 4073 2453 4087 2467
rect 4053 2433 4067 2447
rect 4013 2393 4027 2407
rect 3993 2373 4007 2387
rect 3973 2313 3987 2327
rect 3933 2293 3947 2307
rect 4053 2293 4067 2307
rect 3913 2273 3927 2287
rect 3953 2273 3967 2287
rect 3933 2253 3947 2267
rect 3853 2233 3867 2247
rect 3833 2193 3847 2207
rect 3793 2133 3807 2147
rect 3813 2133 3827 2147
rect 3933 2133 3947 2147
rect 3813 2093 3827 2107
rect 3833 2093 3847 2107
rect 3793 2073 3807 2087
rect 3873 2073 3887 2087
rect 3793 2013 3807 2027
rect 3813 2013 3827 2027
rect 3773 1773 3787 1787
rect 3733 1753 3747 1767
rect 3753 1753 3767 1767
rect 3813 1833 3827 1847
rect 3913 2053 3927 2067
rect 3893 1933 3907 1947
rect 3853 1793 3867 1807
rect 3813 1773 3827 1787
rect 3873 1773 3887 1787
rect 3813 1753 3827 1767
rect 3793 1713 3807 1727
rect 3793 1673 3807 1687
rect 3773 1633 3787 1647
rect 3713 1533 3727 1547
rect 3613 1493 3627 1507
rect 3593 1453 3607 1467
rect 3653 1453 3667 1467
rect 3613 1313 3627 1327
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3593 1273 3607 1287
rect 3613 1273 3627 1287
rect 3633 1273 3647 1287
rect 3613 1233 3627 1247
rect 3573 1113 3587 1127
rect 3593 1113 3607 1127
rect 3533 813 3547 827
rect 3753 1613 3767 1627
rect 3793 1573 3807 1587
rect 3773 1553 3787 1567
rect 3733 1333 3747 1347
rect 3713 1293 3727 1307
rect 3753 1313 3767 1327
rect 3673 1273 3687 1287
rect 3693 1273 3707 1287
rect 3693 1093 3707 1107
rect 3653 973 3667 987
rect 3633 853 3647 867
rect 3713 853 3727 867
rect 3593 813 3607 827
rect 3633 813 3647 827
rect 3513 673 3527 687
rect 3713 793 3727 807
rect 3393 653 3407 667
rect 3453 653 3467 667
rect 3493 653 3507 667
rect 3573 653 3587 667
rect 3413 633 3427 647
rect 3373 613 3387 627
rect 3453 613 3467 627
rect 3533 633 3547 647
rect 3513 613 3527 627
rect 3553 613 3567 627
rect 3673 673 3687 687
rect 3873 1733 3887 1747
rect 3853 1693 3867 1707
rect 3833 1653 3847 1667
rect 4013 2253 4027 2267
rect 4033 2273 4047 2287
rect 3973 2233 3987 2247
rect 3993 2233 4007 2247
rect 4013 2213 4027 2227
rect 4033 2213 4047 2227
rect 3973 2073 3987 2087
rect 3993 1953 4007 1967
rect 3953 1813 3967 1827
rect 3913 1793 3927 1807
rect 3953 1793 3967 1807
rect 3973 1773 3987 1787
rect 4053 2093 4067 2107
rect 4033 2073 4047 2087
rect 4053 2013 4067 2027
rect 4013 1933 4027 1947
rect 4173 2713 4187 2727
rect 4193 2713 4207 2727
rect 4153 2673 4167 2687
rect 4133 2653 4147 2667
rect 4113 2433 4127 2447
rect 4153 2613 4167 2627
rect 4133 2333 4147 2347
rect 4153 2233 4167 2247
rect 4093 2073 4107 2087
rect 4073 1953 4087 1967
rect 4113 1853 4127 1867
rect 3953 1713 3967 1727
rect 3893 1673 3907 1687
rect 3893 1653 3907 1667
rect 3933 1613 3947 1627
rect 3833 1593 3847 1607
rect 3833 1573 3847 1587
rect 3873 1573 3887 1587
rect 3813 1553 3827 1567
rect 3993 1733 4007 1747
rect 4033 1773 4047 1787
rect 4033 1753 4047 1767
rect 4053 1753 4067 1767
rect 4013 1713 4027 1727
rect 3993 1593 4007 1607
rect 4113 1773 4127 1787
rect 4073 1733 4087 1747
rect 4073 1693 4087 1707
rect 4093 1693 4107 1707
rect 4053 1653 4067 1667
rect 4093 1653 4107 1667
rect 4113 1653 4127 1667
rect 4013 1573 4027 1587
rect 3813 1293 3827 1307
rect 3793 1273 3807 1287
rect 3853 1333 3867 1347
rect 3873 1333 3887 1347
rect 3953 1333 3967 1347
rect 3933 1293 3947 1307
rect 3873 1253 3887 1267
rect 4073 1613 4087 1627
rect 4093 1613 4107 1627
rect 4153 1933 4167 1947
rect 4153 1653 4167 1667
rect 4233 2713 4247 2727
rect 4233 2693 4247 2707
rect 4213 2633 4227 2647
rect 4193 2533 4207 2547
rect 4213 2533 4227 2547
rect 4273 2713 4287 2727
rect 4253 2513 4267 2527
rect 4233 2473 4247 2487
rect 4213 2253 4227 2267
rect 4233 2233 4247 2247
rect 4313 2933 4327 2947
rect 4313 2693 4327 2707
rect 4393 3113 4407 3127
rect 4433 3173 4447 3187
rect 4413 3073 4427 3087
rect 4393 3053 4407 3067
rect 4373 2733 4387 2747
rect 4413 3033 4427 3047
rect 4413 3013 4427 3027
rect 4413 2953 4427 2967
rect 4433 2873 4447 2887
rect 4413 2713 4427 2727
rect 4433 2713 4447 2727
rect 4393 2633 4407 2647
rect 4313 2553 4327 2567
rect 4333 2533 4347 2547
rect 4313 2513 4327 2527
rect 4333 2293 4347 2307
rect 4193 2093 4207 2107
rect 4293 2133 4307 2147
rect 4313 2113 4327 2127
rect 4433 2533 4447 2547
rect 4433 2513 4447 2527
rect 4413 2253 4427 2267
rect 4373 2133 4387 2147
rect 4413 2133 4427 2147
rect 4333 2093 4347 2107
rect 4353 2093 4367 2107
rect 4413 2093 4427 2107
rect 4313 2053 4327 2067
rect 4333 2053 4347 2067
rect 4193 1933 4207 1947
rect 4193 1913 4207 1927
rect 4233 1913 4247 1927
rect 4093 1573 4107 1587
rect 4053 1533 4067 1547
rect 4053 1313 4067 1327
rect 4093 1313 4107 1327
rect 4073 1293 4087 1307
rect 4033 1233 4047 1247
rect 3933 1193 3947 1207
rect 4013 1193 4027 1207
rect 3813 1133 3827 1147
rect 3853 1133 3867 1147
rect 3893 1133 3907 1147
rect 3793 813 3807 827
rect 3773 713 3787 727
rect 3673 633 3687 647
rect 3873 1113 3887 1127
rect 3833 1093 3847 1107
rect 3853 1093 3867 1107
rect 3913 1113 3927 1127
rect 3893 1093 3907 1107
rect 3913 973 3927 987
rect 3853 793 3867 807
rect 4013 1113 4027 1127
rect 3973 1093 3987 1107
rect 4033 1093 4047 1107
rect 3953 973 3967 987
rect 3933 853 3947 867
rect 3933 773 3947 787
rect 3833 673 3847 687
rect 3933 673 3947 687
rect 3813 653 3827 667
rect 3813 613 3827 627
rect 3873 633 3887 647
rect 3913 633 3927 647
rect 3893 613 3907 627
rect 3793 533 3807 547
rect 3473 413 3487 427
rect 3613 393 3627 407
rect 3633 393 3647 407
rect 3793 393 3807 407
rect 3113 373 3127 387
rect 3353 373 3367 387
rect 3393 373 3407 387
rect 3473 373 3487 387
rect 3073 353 3087 367
rect 3133 333 3147 347
rect 3173 333 3187 347
rect 3313 353 3327 367
rect 3053 313 3067 327
rect 3093 293 3107 307
rect 3073 213 3087 227
rect 3033 193 3047 207
rect 3033 173 3047 187
rect 3073 153 3087 167
rect 3113 153 3127 167
rect 3233 333 3247 347
rect 3353 353 3367 367
rect 3433 353 3447 367
rect 3193 273 3207 287
rect 3273 253 3287 267
rect 3413 313 3427 327
rect 3453 313 3467 327
rect 3513 333 3527 347
rect 3353 293 3367 307
rect 3493 293 3507 307
rect 3333 233 3347 247
rect 3153 213 3167 227
rect 3193 193 3207 207
rect 3133 133 3147 147
rect 3273 153 3287 167
rect 3233 133 3247 147
rect 3533 313 3547 327
rect 3513 273 3527 287
rect 3393 173 3407 187
rect 3613 333 3627 347
rect 3693 353 3707 367
rect 3593 313 3607 327
rect 3653 313 3667 327
rect 3753 373 3767 387
rect 3773 353 3787 367
rect 3573 293 3587 307
rect 3733 293 3747 307
rect 3573 253 3587 267
rect 3473 153 3487 167
rect 3533 153 3547 167
rect 3733 233 3747 247
rect 3573 153 3587 167
rect 3613 153 3627 167
rect 3693 173 3707 187
rect 3793 173 3807 187
rect 4053 1073 4067 1087
rect 4013 853 4027 867
rect 4033 853 4047 867
rect 3973 833 3987 847
rect 3993 813 4007 827
rect 4073 813 4087 827
rect 4073 773 4087 787
rect 4173 1613 4187 1627
rect 4333 2033 4347 2047
rect 4273 1833 4287 1847
rect 4213 1793 4227 1807
rect 4253 1793 4267 1807
rect 4293 1793 4307 1807
rect 4233 1753 4247 1767
rect 4513 3273 4527 3287
rect 4473 3253 4487 3267
rect 4493 3233 4507 3247
rect 4473 3073 4487 3087
rect 4493 3073 4507 3087
rect 4553 3493 4567 3507
rect 4473 2853 4487 2867
rect 4493 2773 4507 2787
rect 4533 3033 4547 3047
rect 4593 3473 4607 3487
rect 4713 4453 4727 4467
rect 4733 4433 4747 4447
rect 4673 4293 4687 4307
rect 4633 4113 4647 4127
rect 4673 3973 4687 3987
rect 4633 3953 4647 3967
rect 4633 3913 4647 3927
rect 4733 4293 4747 4307
rect 4713 4193 4727 4207
rect 4713 3973 4727 3987
rect 4693 3753 4707 3767
rect 4633 3713 4647 3727
rect 4673 3673 4687 3687
rect 4653 3653 4667 3667
rect 4633 3513 4647 3527
rect 4653 3493 4667 3507
rect 4673 3513 4687 3527
rect 4693 3493 4707 3507
rect 4673 3473 4687 3487
rect 4553 2973 4567 2987
rect 4653 3453 4667 3467
rect 4633 3293 4647 3307
rect 4673 3273 4687 3287
rect 4653 3253 4667 3267
rect 4673 3233 4687 3247
rect 4653 3193 4667 3207
rect 4653 3093 4667 3107
rect 4633 3073 4647 3087
rect 4653 3073 4667 3087
rect 4693 3213 4707 3227
rect 4673 3053 4687 3067
rect 4613 3033 4627 3047
rect 4613 3013 4627 3027
rect 4673 3033 4687 3047
rect 4773 3713 4787 3727
rect 4753 3493 4767 3507
rect 4733 3233 4747 3247
rect 4733 3213 4747 3227
rect 4733 3173 4747 3187
rect 4733 3053 4747 3067
rect 4693 3013 4707 3027
rect 4593 2993 4607 3007
rect 4653 2993 4667 3007
rect 4673 2993 4687 3007
rect 4613 2913 4627 2927
rect 4693 2973 4707 2987
rect 4553 2793 4567 2807
rect 4613 2793 4627 2807
rect 4673 2793 4687 2807
rect 4573 2733 4587 2747
rect 4533 2713 4547 2727
rect 4593 2713 4607 2727
rect 4553 2693 4567 2707
rect 4513 2673 4527 2687
rect 4473 2573 4487 2587
rect 4513 2553 4527 2567
rect 4533 2553 4547 2567
rect 4453 2493 4467 2507
rect 4633 2773 4647 2787
rect 4633 2733 4647 2747
rect 4593 2553 4607 2567
rect 4613 2553 4627 2567
rect 4553 2513 4567 2527
rect 4573 2513 4587 2527
rect 4673 2733 4687 2747
rect 4653 2713 4667 2727
rect 4693 2693 4707 2707
rect 4613 2513 4627 2527
rect 4633 2513 4647 2527
rect 4693 2513 4707 2527
rect 4493 2473 4507 2487
rect 4653 2493 4667 2507
rect 4613 2473 4627 2487
rect 4453 2253 4467 2267
rect 4573 2333 4587 2347
rect 4693 2473 4707 2487
rect 4573 2313 4587 2327
rect 4533 2293 4547 2307
rect 4613 2273 4627 2287
rect 4593 2253 4607 2267
rect 4553 2173 4567 2187
rect 4693 2313 4707 2327
rect 4653 2293 4667 2307
rect 4673 2273 4687 2287
rect 4673 2253 4687 2267
rect 4533 2153 4547 2167
rect 4593 2153 4607 2167
rect 4533 2133 4547 2147
rect 4473 2113 4487 2127
rect 4493 2093 4507 2107
rect 4373 2053 4387 2067
rect 4513 2073 4527 2087
rect 4493 2053 4507 2067
rect 4353 1793 4367 1807
rect 4333 1773 4347 1787
rect 4233 1733 4247 1747
rect 4213 1693 4227 1707
rect 4273 1693 4287 1707
rect 4293 1673 4307 1687
rect 4273 1653 4287 1667
rect 4253 1613 4267 1627
rect 4213 1573 4227 1587
rect 4253 1573 4267 1587
rect 4133 1533 4147 1547
rect 4193 1533 4207 1547
rect 4173 1393 4187 1407
rect 4173 1373 4187 1387
rect 4133 1353 4147 1367
rect 4153 1313 4167 1327
rect 4133 1133 4147 1147
rect 4173 1133 4187 1147
rect 4253 1533 4267 1547
rect 4213 1493 4227 1507
rect 4413 1773 4427 1787
rect 4333 1693 4347 1707
rect 4313 1653 4327 1667
rect 4393 1753 4407 1767
rect 4393 1733 4407 1747
rect 4333 1613 4347 1627
rect 4353 1613 4367 1627
rect 4353 1573 4367 1587
rect 4373 1593 4387 1607
rect 4313 1553 4327 1567
rect 4353 1553 4367 1567
rect 4253 1413 4267 1427
rect 4293 1413 4307 1427
rect 4213 1353 4227 1367
rect 4193 1073 4207 1087
rect 4113 793 4127 807
rect 4033 673 4047 687
rect 4013 653 4027 667
rect 3953 633 3967 647
rect 3973 613 3987 627
rect 3993 593 4007 607
rect 3913 573 3927 587
rect 3993 533 4007 547
rect 3893 413 3907 427
rect 3833 353 3847 367
rect 3853 333 3867 347
rect 3873 273 3887 287
rect 3933 293 3947 307
rect 3973 293 3987 307
rect 3913 253 3927 267
rect 3833 173 3847 187
rect 3813 153 3827 167
rect 3973 253 3987 267
rect 3953 213 3967 227
rect 3873 153 3887 167
rect 3893 153 3907 167
rect 3793 133 3807 147
rect 3913 113 3927 127
rect 4033 633 4047 647
rect 4033 593 4047 607
rect 4093 633 4107 647
rect 4093 573 4107 587
rect 4073 353 4087 367
rect 4033 313 4047 327
rect 4073 333 4087 347
rect 4113 333 4127 347
rect 4153 793 4167 807
rect 4173 793 4187 807
rect 4153 633 4167 647
rect 4293 1393 4307 1407
rect 4373 1513 4387 1527
rect 4273 1173 4287 1187
rect 4333 1313 4347 1327
rect 4413 1673 4427 1687
rect 4453 1793 4467 1807
rect 4513 1833 4527 1847
rect 4493 1773 4507 1787
rect 4453 1713 4467 1727
rect 4413 1653 4427 1667
rect 4433 1653 4447 1667
rect 4433 1573 4447 1587
rect 4473 1693 4487 1707
rect 4553 2073 4567 2087
rect 4553 1833 4567 1847
rect 4573 1773 4587 1787
rect 4633 2133 4647 2147
rect 4593 1733 4607 1747
rect 4733 3013 4747 3027
rect 4773 3073 4787 3087
rect 4773 3053 4787 3067
rect 4773 2913 4787 2927
rect 4753 2733 4767 2747
rect 4773 2333 4787 2347
rect 4733 2253 4747 2267
rect 4653 1813 4667 1827
rect 4733 1813 4747 1827
rect 4673 1773 4687 1787
rect 4653 1713 4667 1727
rect 4653 1673 4667 1687
rect 4533 1653 4547 1667
rect 4513 1613 4527 1627
rect 4513 1593 4527 1607
rect 4493 1573 4507 1587
rect 4453 1553 4467 1567
rect 4473 1553 4487 1567
rect 4393 1373 4407 1387
rect 4473 1353 4487 1367
rect 4393 1313 4407 1327
rect 4373 1293 4387 1307
rect 4413 1293 4427 1307
rect 4433 1313 4447 1327
rect 4573 1613 4587 1627
rect 4593 1593 4607 1607
rect 4613 1573 4627 1587
rect 4633 1593 4647 1607
rect 4673 1593 4687 1607
rect 4713 1593 4727 1607
rect 4753 1593 4767 1607
rect 4773 1593 4787 1607
rect 4633 1513 4647 1527
rect 4693 1553 4707 1567
rect 4713 1573 4727 1587
rect 4733 1553 4747 1567
rect 4633 1353 4647 1367
rect 4673 1353 4687 1367
rect 4693 1353 4707 1367
rect 4453 1253 4467 1267
rect 4433 1153 4447 1167
rect 4393 1133 4407 1147
rect 4293 1113 4307 1127
rect 4333 1113 4347 1127
rect 4353 1113 4367 1127
rect 4273 1073 4287 1087
rect 4293 1093 4307 1107
rect 4373 1093 4387 1107
rect 4413 1093 4427 1107
rect 4493 1293 4507 1307
rect 4533 1313 4547 1327
rect 4553 1293 4567 1307
rect 4513 1273 4527 1287
rect 4673 1313 4687 1327
rect 4573 1273 4587 1287
rect 4593 1253 4607 1267
rect 4573 1153 4587 1167
rect 4553 1133 4567 1147
rect 4653 1273 4667 1287
rect 4433 1073 4447 1087
rect 4253 813 4267 827
rect 4313 813 4327 827
rect 4193 753 4207 767
rect 4213 713 4227 727
rect 4233 613 4247 627
rect 4213 593 4227 607
rect 4253 593 4267 607
rect 4273 613 4287 627
rect 4493 1113 4507 1127
rect 4473 1073 4487 1087
rect 4493 1093 4507 1107
rect 4553 1093 4567 1107
rect 4633 1113 4647 1127
rect 4593 1093 4607 1107
rect 4733 1333 4747 1347
rect 4773 1573 4787 1587
rect 4773 1353 4787 1367
rect 4713 1313 4727 1327
rect 4753 1313 4767 1327
rect 4773 1313 4787 1327
rect 4673 1113 4687 1127
rect 4693 1113 4707 1127
rect 4553 1073 4567 1087
rect 4513 1033 4527 1047
rect 4493 913 4507 927
rect 4453 813 4467 827
rect 4413 793 4427 807
rect 4373 773 4387 787
rect 4653 1073 4667 1087
rect 4673 1053 4687 1067
rect 4613 913 4627 927
rect 4653 913 4667 927
rect 4553 893 4567 907
rect 4613 873 4627 887
rect 4693 1033 4707 1047
rect 4673 853 4687 867
rect 4453 753 4467 767
rect 4393 673 4407 687
rect 4353 613 4367 627
rect 4493 673 4507 687
rect 4433 613 4447 627
rect 4133 313 4147 327
rect 4113 293 4127 307
rect 4033 253 4047 267
rect 3993 173 4007 187
rect 4013 173 4027 187
rect 3993 153 4007 167
rect 4073 153 4087 167
rect 4473 513 4487 527
rect 4633 813 4647 827
rect 4753 1133 4767 1147
rect 4733 1113 4747 1127
rect 4753 913 4767 927
rect 4753 893 4767 907
rect 4733 873 4747 887
rect 4633 793 4647 807
rect 4673 793 4687 807
rect 4693 773 4707 787
rect 4293 413 4307 427
rect 4473 413 4487 427
rect 4533 413 4547 427
rect 4273 393 4287 407
rect 4353 393 4367 407
rect 4253 333 4267 347
rect 4193 273 4207 287
rect 4173 173 4187 187
rect 4193 173 4207 187
rect 4053 133 4067 147
rect 4313 373 4327 387
rect 4333 353 4347 367
rect 4373 373 4387 387
rect 4393 333 4407 347
rect 4433 353 4447 367
rect 4493 353 4507 367
rect 4473 313 4487 327
rect 4413 293 4427 307
rect 4373 213 4387 227
rect 4333 173 4347 187
rect 4213 153 4227 167
rect 4253 133 4267 147
rect 4293 133 4307 147
rect 3973 113 3987 127
rect 4413 173 4427 187
rect 4453 173 4467 187
rect 4653 633 4667 647
rect 4673 633 4687 647
rect 4513 193 4527 207
rect 4493 173 4507 187
rect 4513 173 4527 187
rect 4613 173 4627 187
rect 4713 633 4727 647
rect 4693 513 4707 527
rect 4673 293 4687 307
rect 4433 133 4447 147
rect 4473 153 4487 167
rect 4533 153 4547 167
rect 4573 133 4587 147
rect 4653 133 4667 147
rect 4693 113 4707 127
rect 4753 133 4767 147
rect 4433 93 4447 107
rect 4733 93 4747 107
rect 1973 13 1987 27
rect 2113 13 2127 27
rect 2153 13 2167 27
<< metal3 >>
rect 4067 4576 4113 4584
rect 4147 4576 4233 4584
rect 4327 4576 4353 4584
rect 1247 4556 1533 4564
rect 4047 4556 4153 4564
rect 127 4536 193 4544
rect 907 4536 1293 4544
rect 1467 4536 1633 4544
rect 2287 4536 2333 4544
rect 3347 4536 3433 4544
rect 3967 4536 4193 4544
rect 47 4516 493 4524
rect 727 4516 1433 4524
rect 1447 4516 1613 4524
rect 1627 4516 1693 4524
rect 1707 4516 1813 4524
rect 1967 4516 2013 4524
rect 2067 4516 2293 4524
rect 3027 4516 3053 4524
rect 3107 4516 3173 4524
rect 3247 4516 3493 4524
rect 3987 4516 4613 4524
rect 87 4496 173 4504
rect 387 4496 433 4504
rect 567 4496 644 4504
rect 187 4476 213 4484
rect 407 4476 444 4484
rect 107 4456 153 4464
rect 167 4456 233 4464
rect 267 4456 313 4464
rect 367 4456 413 4464
rect 436 4464 444 4476
rect 487 4476 604 4484
rect 436 4456 453 4464
rect 467 4456 493 4464
rect 287 4436 373 4444
rect 496 4436 513 4444
rect 527 4436 533 4444
rect 107 4416 153 4424
rect 176 4424 184 4433
rect 176 4416 193 4424
rect 596 4424 604 4476
rect 636 4484 644 4496
rect 667 4496 1053 4504
rect 1087 4496 1113 4504
rect 1147 4496 1273 4504
rect 1327 4496 1353 4504
rect 1376 4496 1453 4504
rect 636 4476 753 4484
rect 787 4476 833 4484
rect 867 4476 984 4484
rect 616 4447 624 4473
rect 707 4456 753 4464
rect 867 4456 933 4464
rect 976 4464 984 4476
rect 1007 4476 1104 4484
rect 1096 4467 1104 4476
rect 1167 4476 1173 4484
rect 1187 4476 1333 4484
rect 1376 4484 1384 4496
rect 1567 4496 1773 4504
rect 1896 4496 1913 4504
rect 1356 4476 1384 4484
rect 976 4456 1033 4464
rect 1047 4456 1084 4464
rect 676 4444 684 4453
rect 667 4436 684 4444
rect 596 4416 633 4424
rect 796 4424 804 4453
rect 816 4427 824 4453
rect 847 4436 864 4444
rect 856 4427 864 4436
rect 887 4436 904 4444
rect 727 4416 804 4424
rect 67 4396 113 4404
rect 127 4396 173 4404
rect 347 4396 693 4404
rect 896 4404 904 4436
rect 967 4436 1013 4444
rect 1076 4444 1084 4456
rect 1107 4456 1193 4464
rect 1356 4464 1364 4476
rect 1407 4476 1484 4484
rect 1287 4456 1364 4464
rect 1476 4464 1484 4476
rect 1507 4476 1573 4484
rect 1896 4484 1904 4496
rect 1927 4496 2173 4504
rect 2196 4496 2393 4504
rect 1587 4476 1904 4484
rect 2196 4484 2204 4496
rect 2407 4496 2473 4504
rect 2947 4496 2993 4504
rect 3007 4496 3113 4504
rect 3127 4496 3133 4504
rect 3187 4496 3413 4504
rect 3427 4496 3464 4504
rect 2007 4476 2204 4484
rect 2227 4476 2324 4484
rect 2316 4467 2324 4476
rect 2516 4484 2524 4493
rect 3456 4487 3464 4496
rect 3647 4496 4133 4504
rect 4167 4496 4333 4504
rect 2447 4476 2524 4484
rect 2667 4476 2793 4484
rect 3016 4476 3144 4484
rect 1476 4456 1553 4464
rect 1607 4456 1653 4464
rect 1907 4456 2013 4464
rect 2147 4456 2193 4464
rect 1076 4436 1133 4444
rect 1376 4444 1384 4453
rect 1267 4436 1384 4444
rect 1527 4436 1693 4444
rect 1847 4436 1973 4444
rect 2267 4436 2353 4444
rect 2376 4444 2384 4473
rect 2616 4464 2624 4473
rect 2467 4456 2624 4464
rect 2727 4456 2973 4464
rect 3016 4464 3024 4476
rect 2987 4456 3024 4464
rect 3087 4456 3113 4464
rect 3136 4464 3144 4476
rect 3287 4476 3353 4484
rect 3367 4476 3373 4484
rect 3587 4476 3713 4484
rect 4127 4476 4273 4484
rect 4327 4476 4513 4484
rect 3136 4456 3253 4464
rect 3267 4456 3293 4464
rect 3407 4456 3693 4464
rect 3747 4456 3793 4464
rect 4247 4456 4293 4464
rect 4687 4456 4713 4464
rect 2376 4436 2493 4444
rect 2547 4436 2673 4444
rect 3036 4444 3044 4453
rect 3036 4436 3073 4444
rect 3667 4436 3773 4444
rect 3787 4436 4093 4444
rect 4187 4436 4293 4444
rect 4627 4436 4733 4444
rect 927 4416 1093 4424
rect 1187 4416 1284 4424
rect 896 4396 1044 4404
rect 667 4376 733 4384
rect 1036 4384 1044 4396
rect 1067 4396 1253 4404
rect 1276 4404 1284 4416
rect 1367 4416 1593 4424
rect 1607 4416 2433 4424
rect 2587 4416 2633 4424
rect 3027 4416 3193 4424
rect 3807 4416 4053 4424
rect 1276 4396 1413 4404
rect 1567 4396 1753 4404
rect 1767 4396 2033 4404
rect 2427 4396 4033 4404
rect 4207 4396 4393 4404
rect 1036 4376 1213 4384
rect 2467 4376 3953 4384
rect 147 4356 553 4364
rect 567 4356 593 4364
rect 607 4356 813 4364
rect 827 4356 913 4364
rect 967 4356 1073 4364
rect 1087 4356 1153 4364
rect 467 4316 573 4324
rect 1807 4316 1893 4324
rect 1907 4316 1933 4324
rect 1947 4316 2093 4324
rect 4047 4296 4093 4304
rect 4107 4296 4133 4304
rect 4687 4296 4733 4304
rect 367 4276 413 4284
rect 2127 4276 3193 4284
rect 1687 4256 2004 4264
rect 47 4236 93 4244
rect 1407 4236 1484 4244
rect 1476 4227 1484 4236
rect 1567 4236 1793 4244
rect 1807 4236 1933 4244
rect 87 4216 124 4224
rect 96 4184 104 4193
rect 87 4176 104 4184
rect 116 4167 124 4216
rect 167 4216 184 4224
rect 176 4204 184 4216
rect 227 4216 264 4224
rect 147 4196 164 4204
rect 176 4196 233 4204
rect 156 4184 164 4196
rect 256 4204 264 4216
rect 327 4216 504 4224
rect 256 4196 284 4204
rect 156 4176 253 4184
rect 276 4184 284 4196
rect 316 4196 413 4204
rect 276 4176 293 4184
rect 316 4167 324 4196
rect 427 4196 473 4204
rect 496 4204 504 4216
rect 667 4216 724 4224
rect 496 4196 513 4204
rect 716 4204 724 4216
rect 807 4216 913 4224
rect 1067 4216 1113 4224
rect 1307 4216 1433 4224
rect 1447 4216 1464 4224
rect 1456 4207 1464 4216
rect 1927 4216 1973 4224
rect 716 4196 773 4204
rect 1247 4196 1313 4204
rect 1467 4196 1553 4204
rect 1747 4196 1813 4204
rect 367 4176 393 4184
rect 696 4184 704 4193
rect 507 4176 813 4184
rect 867 4176 893 4184
rect 956 4184 964 4193
rect 956 4176 1093 4184
rect 1247 4176 1273 4184
rect 1347 4176 1393 4184
rect 1836 4184 1844 4213
rect 1767 4176 1844 4184
rect 567 4156 673 4164
rect 707 4156 713 4164
rect 727 4156 753 4164
rect 887 4156 933 4164
rect 1507 4156 1673 4164
rect 1876 4164 1884 4213
rect 1996 4204 2004 4256
rect 3127 4256 3253 4264
rect 2687 4236 3273 4244
rect 3407 4236 3493 4244
rect 3667 4236 3713 4244
rect 3727 4236 4193 4244
rect 4227 4236 4553 4244
rect 2027 4216 2104 4224
rect 2096 4207 2104 4216
rect 2927 4216 3093 4224
rect 3327 4216 3613 4224
rect 3627 4216 3673 4224
rect 3947 4216 4133 4224
rect 4296 4216 4353 4224
rect 1936 4196 2004 4204
rect 1896 4184 1904 4193
rect 1936 4187 1944 4196
rect 2507 4196 2864 4204
rect 1896 4176 1924 4184
rect 1687 4156 1893 4164
rect 1916 4164 1924 4176
rect 2367 4176 2553 4184
rect 2607 4176 2633 4184
rect 2856 4184 2864 4196
rect 2887 4196 3013 4204
rect 3067 4196 3113 4204
rect 3236 4204 3244 4213
rect 3236 4196 3293 4204
rect 3827 4196 3833 4204
rect 3847 4196 3944 4204
rect 2856 4176 2933 4184
rect 3016 4184 3024 4193
rect 2987 4176 3024 4184
rect 3227 4176 3493 4184
rect 3627 4176 3773 4184
rect 3887 4176 3913 4184
rect 3936 4184 3944 4196
rect 3936 4176 4053 4184
rect 1916 4156 1973 4164
rect 2527 4156 2553 4164
rect 2607 4156 2853 4164
rect 2967 4156 3073 4164
rect 3087 4156 3093 4164
rect 3267 4156 3333 4164
rect 3387 4156 3433 4164
rect 3667 4156 3733 4164
rect 3787 4156 4013 4164
rect 4176 4164 4184 4193
rect 4296 4184 4304 4216
rect 4327 4196 4433 4204
rect 4487 4196 4713 4204
rect 4287 4176 4304 4184
rect 4387 4176 4513 4184
rect 4087 4156 4184 4164
rect 4207 4156 4333 4164
rect 4347 4156 4453 4164
rect 67 4136 293 4144
rect 607 4136 773 4144
rect 907 4136 1033 4144
rect 1047 4136 1133 4144
rect 1207 4136 1453 4144
rect 1867 4136 2073 4144
rect 2927 4136 2953 4144
rect 2967 4136 2993 4144
rect 3927 4136 4493 4144
rect 4507 4136 4513 4144
rect 4527 4136 4593 4144
rect 187 4116 373 4124
rect 527 4116 593 4124
rect 1087 4116 1333 4124
rect 1427 4116 1713 4124
rect 1727 4116 2133 4124
rect 2147 4116 2173 4124
rect 2767 4116 3033 4124
rect 3167 4116 4373 4124
rect 4427 4116 4633 4124
rect 167 4096 433 4104
rect 1367 4096 1413 4104
rect 1627 4096 1653 4104
rect 1667 4096 1713 4104
rect 2007 4096 2073 4104
rect 2087 4096 2313 4104
rect 3567 4096 3693 4104
rect 4047 4096 4213 4104
rect 4247 4096 4293 4104
rect 167 4076 273 4084
rect 287 4076 333 4084
rect 1547 4076 1873 4084
rect 2287 4076 2713 4084
rect 2727 4076 2813 4084
rect 2827 4076 3533 4084
rect 3547 4076 3653 4084
rect 3667 4076 3873 4084
rect 4287 4076 4333 4084
rect 207 4056 293 4064
rect 667 4056 793 4064
rect 807 4056 1073 4064
rect 1827 4056 2253 4064
rect 3367 4056 4033 4064
rect 4047 4056 4073 4064
rect 4107 4056 4133 4064
rect 4147 4056 4193 4064
rect 67 4036 373 4044
rect 427 4036 853 4044
rect 867 4036 933 4044
rect 967 4036 1213 4044
rect 1227 4036 1373 4044
rect 1807 4036 1933 4044
rect 2067 4036 2273 4044
rect 2287 4036 2373 4044
rect 2747 4036 2993 4044
rect 3247 4036 3673 4044
rect 3867 4036 3933 4044
rect 3947 4036 4093 4044
rect 87 4016 213 4024
rect 347 4016 493 4024
rect 507 4016 644 4024
rect 447 3996 513 4004
rect 536 3996 613 4004
rect 267 3976 273 3984
rect 536 3984 544 3996
rect 636 3987 644 4016
rect 727 4016 1233 4024
rect 1247 4016 1353 4024
rect 1367 4016 1433 4024
rect 1487 4016 1544 4024
rect 736 3996 773 4004
rect 287 3976 544 3984
rect 567 3976 624 3984
rect 47 3956 193 3964
rect 276 3964 284 3973
rect 276 3956 353 3964
rect 616 3964 624 3976
rect 676 3964 684 3973
rect 616 3956 684 3964
rect 147 3936 453 3944
rect 467 3936 573 3944
rect 736 3944 744 3996
rect 1007 3996 1013 4004
rect 1407 3996 1513 4004
rect 767 3976 813 3984
rect 956 3976 973 3984
rect 756 3947 764 3973
rect 787 3956 833 3964
rect 667 3936 744 3944
rect 836 3944 844 3953
rect 836 3936 873 3944
rect 956 3944 964 3976
rect 996 3964 1004 3993
rect 1047 3976 1133 3984
rect 1307 3976 1333 3984
rect 987 3956 1004 3964
rect 1107 3956 1193 3964
rect 1407 3956 1453 3964
rect 1536 3964 1544 4016
rect 1667 4016 1813 4024
rect 1927 4016 1953 4024
rect 2407 4016 2433 4024
rect 2587 4016 3053 4024
rect 3087 4016 3213 4024
rect 3227 4016 3273 4024
rect 3287 4016 3313 4024
rect 3347 4016 3453 4024
rect 3487 4016 3753 4024
rect 3836 4016 3913 4024
rect 1607 3996 1633 4004
rect 1687 3996 1693 4004
rect 1707 3996 1753 4004
rect 2287 3996 2353 4004
rect 3107 3996 3244 4004
rect 1507 3956 1544 3964
rect 956 3936 1033 3944
rect 1427 3936 1473 3944
rect 1487 3936 1533 3944
rect 1776 3944 1784 3993
rect 1836 3967 1844 3993
rect 1927 3976 1973 3984
rect 2107 3976 2153 3984
rect 2227 3976 2293 3984
rect 2776 3984 2784 3993
rect 2627 3976 2784 3984
rect 2927 3976 2973 3984
rect 3027 3976 3153 3984
rect 3236 3984 3244 3996
rect 3387 3996 3413 4004
rect 3707 3996 3813 4004
rect 3236 3976 3253 3984
rect 3356 3967 3364 3993
rect 3436 3984 3444 3993
rect 3836 3987 3844 4016
rect 4027 4016 4153 4024
rect 3856 3996 3893 4004
rect 3856 3987 3864 3996
rect 4007 3996 4053 4004
rect 4127 3996 4184 4004
rect 4176 3987 4184 3996
rect 4207 3996 4273 4004
rect 4307 3996 4553 4004
rect 3376 3976 3513 3984
rect 3376 3967 3384 3976
rect 4227 3976 4313 3984
rect 4427 3976 4673 3984
rect 4687 3976 4713 3984
rect 1867 3956 1993 3964
rect 2687 3956 2773 3964
rect 2947 3956 3133 3964
rect 3687 3956 3973 3964
rect 4647 3956 4824 3964
rect 1776 3936 1813 3944
rect 3187 3936 3573 3944
rect 3587 3936 3853 3944
rect 267 3916 433 3924
rect 447 3916 533 3924
rect 707 3916 853 3924
rect 2387 3916 3633 3924
rect 3827 3916 3873 3924
rect 3887 3916 4633 3924
rect 67 3896 313 3904
rect 327 3896 393 3904
rect 547 3896 593 3904
rect 1127 3896 1233 3904
rect 1247 3896 1273 3904
rect 2487 3896 3773 3904
rect 167 3876 173 3884
rect 187 3876 373 3884
rect 1347 3856 1513 3864
rect 1527 3856 1573 3864
rect 4247 3856 4293 3864
rect 3687 3836 4053 3844
rect 4067 3836 4313 3844
rect 887 3796 1033 3804
rect 1047 3796 1173 3804
rect 847 3776 953 3784
rect 427 3756 593 3764
rect 647 3756 993 3764
rect 916 3747 924 3756
rect 1427 3756 1633 3764
rect 1907 3756 1953 3764
rect 3167 3756 3513 3764
rect 3527 3756 3613 3764
rect 4507 3756 4533 3764
rect 4547 3756 4693 3764
rect 407 3736 513 3744
rect 676 3736 844 3744
rect 56 3687 64 3713
rect 76 3707 84 3733
rect 116 3687 124 3713
rect 136 3704 144 3733
rect 167 3716 213 3724
rect 367 3716 493 3724
rect 136 3696 153 3704
rect 296 3704 304 3713
rect 236 3696 304 3704
rect 336 3704 344 3713
rect 516 3707 524 3733
rect 676 3724 684 3736
rect 587 3716 684 3724
rect 747 3716 793 3724
rect 836 3724 844 3736
rect 956 3736 1024 3744
rect 956 3724 964 3736
rect 836 3716 964 3724
rect 1016 3724 1024 3736
rect 1047 3736 1073 3744
rect 1127 3736 1373 3744
rect 1387 3736 1573 3744
rect 1987 3736 2153 3744
rect 2347 3736 2473 3744
rect 3287 3736 3393 3744
rect 3547 3736 3573 3744
rect 4216 3736 4253 3744
rect 1016 3716 1053 3724
rect 1107 3716 1193 3724
rect 1287 3716 1353 3724
rect 1447 3716 1493 3724
rect 1547 3716 1593 3724
rect 1936 3724 1944 3733
rect 1936 3716 2053 3724
rect 2327 3716 2633 3724
rect 3227 3716 3273 3724
rect 3307 3716 3313 3724
rect 3347 3716 3444 3724
rect 336 3696 353 3704
rect 236 3687 244 3696
rect 547 3696 573 3704
rect 267 3676 313 3684
rect 327 3676 413 3684
rect 676 3684 684 3693
rect 696 3687 704 3713
rect 767 3696 933 3704
rect 976 3704 984 3713
rect 976 3696 1013 3704
rect 1067 3696 1133 3704
rect 1487 3696 1513 3704
rect 1676 3704 1684 3713
rect 1567 3696 1684 3704
rect 1707 3696 1713 3704
rect 1727 3696 1733 3704
rect 1756 3687 1764 3713
rect 1787 3696 1813 3704
rect 1827 3696 1953 3704
rect 2147 3696 2373 3704
rect 2507 3696 2533 3704
rect 2547 3696 2613 3704
rect 2676 3687 2684 3713
rect 2727 3696 2873 3704
rect 2976 3704 2984 3713
rect 2927 3696 2984 3704
rect 3156 3704 3164 3713
rect 3156 3696 3253 3704
rect 3316 3704 3324 3713
rect 3316 3696 3344 3704
rect 427 3676 684 3684
rect 847 3676 913 3684
rect 947 3676 973 3684
rect 1087 3676 1173 3684
rect 1227 3676 1253 3684
rect 1407 3676 1413 3684
rect 1427 3676 1453 3684
rect 1587 3676 1613 3684
rect 1627 3676 1653 3684
rect 1887 3676 1913 3684
rect 1967 3676 1993 3684
rect 2467 3676 2653 3684
rect 2767 3676 2793 3684
rect 2907 3676 2953 3684
rect 3087 3676 3193 3684
rect 3336 3684 3344 3696
rect 3436 3687 3444 3716
rect 3907 3716 4193 3724
rect 3716 3704 3724 3713
rect 3567 3696 3724 3704
rect 3747 3696 3873 3704
rect 4216 3704 4224 3736
rect 4247 3716 4273 3724
rect 4647 3716 4773 3724
rect 4196 3696 4224 3704
rect 4196 3687 4204 3696
rect 4267 3696 4433 3704
rect 4816 3704 4824 3724
rect 4796 3696 4824 3704
rect 3336 3676 3373 3684
rect 3707 3676 3773 3684
rect 3807 3676 4073 3684
rect 4796 3684 4804 3696
rect 4687 3676 4804 3684
rect 87 3656 133 3664
rect 187 3656 373 3664
rect 527 3656 933 3664
rect 1267 3656 1553 3664
rect 1847 3656 2393 3664
rect 2607 3656 2753 3664
rect 2967 3656 3113 3664
rect 3127 3656 3353 3664
rect 3467 3656 3813 3664
rect 4127 3656 4213 3664
rect 4816 3664 4824 3684
rect 4667 3656 4824 3664
rect 67 3636 93 3644
rect 247 3636 313 3644
rect 447 3636 453 3644
rect 467 3636 793 3644
rect 1087 3636 1373 3644
rect 1387 3636 1633 3644
rect 1647 3636 1913 3644
rect 2827 3636 2993 3644
rect 3007 3636 3133 3644
rect 3407 3636 3633 3644
rect 4187 3636 4293 3644
rect 47 3616 93 3624
rect 127 3616 373 3624
rect 387 3616 693 3624
rect 767 3616 1133 3624
rect 1147 3616 1573 3624
rect 1947 3616 2373 3624
rect 2787 3616 2913 3624
rect 3307 3616 3413 3624
rect 3427 3616 3433 3624
rect 4167 3616 4273 3624
rect 4327 3616 4413 3624
rect 127 3596 644 3604
rect 347 3576 353 3584
rect 367 3576 533 3584
rect 547 3576 593 3584
rect 636 3584 644 3596
rect 667 3596 1073 3604
rect 1107 3596 1533 3604
rect 2007 3596 2153 3604
rect 2167 3596 2313 3604
rect 3067 3596 3493 3604
rect 3507 3596 3593 3604
rect 3827 3596 4093 3604
rect 4187 3596 4353 3604
rect 4387 3596 4413 3604
rect 636 3576 993 3584
rect 1127 3576 1153 3584
rect 2187 3576 2493 3584
rect 3187 3576 3653 3584
rect 3927 3576 4053 3584
rect -24 3544 -16 3564
rect 687 3556 733 3564
rect 987 3556 1273 3564
rect 1607 3556 2173 3564
rect 2307 3556 2433 3564
rect 2587 3556 2713 3564
rect 3227 3556 3273 3564
rect 3367 3556 3393 3564
rect 3487 3556 3533 3564
rect 3547 3556 3573 3564
rect 3587 3556 3673 3564
rect 4047 3556 4153 3564
rect -44 3536 -16 3544
rect -44 3444 -36 3536
rect 187 3536 513 3544
rect 576 3536 753 3544
rect -24 3504 -16 3524
rect 487 3516 553 3524
rect -24 3496 373 3504
rect 447 3496 493 3504
rect 576 3504 584 3536
rect 847 3536 873 3544
rect 1027 3536 1053 3544
rect 1107 3536 1233 3544
rect 1396 3536 1684 3544
rect 1396 3524 1404 3536
rect 1676 3527 1684 3536
rect 1707 3536 1793 3544
rect 1847 3536 2113 3544
rect 2387 3536 2433 3544
rect 2547 3536 3033 3544
rect 3167 3536 3213 3544
rect 3247 3536 3313 3544
rect 3327 3536 3333 3544
rect 3356 3536 3413 3544
rect 1007 3516 1404 3524
rect 1427 3516 1553 3524
rect 1727 3516 1793 3524
rect 2127 3516 2153 3524
rect 2167 3516 2233 3524
rect 2687 3516 2813 3524
rect 2827 3516 2833 3524
rect 2847 3516 2933 3524
rect 2947 3516 3064 3524
rect 547 3496 584 3504
rect -24 3476 13 3484
rect 87 3476 113 3484
rect 656 3484 664 3513
rect 836 3504 844 3513
rect 836 3496 873 3504
rect 907 3496 1013 3504
rect 1047 3496 1113 3504
rect 1167 3496 1233 3504
rect 1327 3496 1433 3504
rect 1767 3496 1853 3504
rect 2007 3496 2124 3504
rect 567 3476 664 3484
rect 696 3467 704 3493
rect 2116 3487 2124 3496
rect 2267 3496 2333 3504
rect 2407 3496 2693 3504
rect 2747 3496 2873 3504
rect 3056 3504 3064 3516
rect 3087 3516 3133 3524
rect 3187 3516 3253 3524
rect 3356 3524 3364 3536
rect 3447 3536 3464 3544
rect 3336 3516 3364 3524
rect 3456 3524 3464 3536
rect 3487 3536 3513 3544
rect 3556 3536 3653 3544
rect 3456 3516 3504 3524
rect 3056 3496 3193 3504
rect 3336 3504 3344 3516
rect 3247 3496 3344 3504
rect 3407 3496 3433 3504
rect 3496 3487 3504 3516
rect 3556 3507 3564 3536
rect 3767 3536 3913 3544
rect 3967 3536 4033 3544
rect 3627 3516 3804 3524
rect 3796 3507 3804 3516
rect 3867 3516 3953 3524
rect 4067 3516 4293 3524
rect 4307 3516 4393 3524
rect 4487 3516 4633 3524
rect 3727 3496 3753 3504
rect 4407 3496 4453 3504
rect 4567 3496 4653 3504
rect 4676 3487 4684 3513
rect 4707 3496 4753 3504
rect 1007 3476 1033 3484
rect 1107 3476 1193 3484
rect 1267 3476 1293 3484
rect 1347 3476 1373 3484
rect 1607 3476 1673 3484
rect 1687 3476 1893 3484
rect 1927 3476 1953 3484
rect 1967 3476 1973 3484
rect 2907 3476 2953 3484
rect 3187 3476 3293 3484
rect 3567 3476 3693 3484
rect 3707 3476 4593 3484
rect 387 3456 413 3464
rect 427 3456 673 3464
rect 796 3456 1733 3464
rect -44 3436 93 3444
rect 796 3444 804 3456
rect 1767 3456 1813 3464
rect 2027 3456 2093 3464
rect 3007 3456 3233 3464
rect 3787 3456 3833 3464
rect 3847 3456 3893 3464
rect 3947 3456 4013 3464
rect 4027 3456 4333 3464
rect 4367 3456 4653 3464
rect 307 3436 804 3444
rect 827 3436 1073 3444
rect 1867 3436 1893 3444
rect 3847 3436 4073 3444
rect 27 3416 1253 3424
rect 1687 3416 2093 3424
rect 2767 3416 4153 3424
rect 4167 3416 4213 3424
rect 27 3396 293 3404
rect 627 3396 853 3404
rect 947 3396 1013 3404
rect 1227 3396 1473 3404
rect 1487 3396 1713 3404
rect 1727 3396 1773 3404
rect 3307 3396 3873 3404
rect 727 3376 753 3384
rect 767 3376 1004 3384
rect 267 3356 533 3364
rect 687 3356 733 3364
rect 927 3356 973 3364
rect 996 3364 1004 3376
rect 1107 3376 1673 3384
rect 1807 3376 1973 3384
rect 996 3356 1373 3364
rect 1396 3356 1713 3364
rect 267 3336 633 3344
rect 787 3336 1093 3344
rect 1396 3344 1404 3356
rect 1747 3356 1933 3364
rect 2367 3356 2513 3364
rect 1147 3336 1404 3344
rect 1447 3336 2153 3344
rect 3487 3336 3533 3344
rect 327 3316 393 3324
rect 467 3316 513 3324
rect 527 3316 1213 3324
rect 1647 3316 2133 3324
rect 3167 3316 3473 3324
rect 3607 3316 3773 3324
rect 4087 3316 4493 3324
rect 467 3296 553 3304
rect 607 3296 824 3304
rect 47 3276 293 3284
rect 347 3276 393 3284
rect 407 3276 793 3284
rect 816 3284 824 3296
rect 847 3296 1133 3304
rect 1187 3296 1833 3304
rect 2287 3296 2333 3304
rect 2347 3296 2393 3304
rect 3287 3296 3573 3304
rect 3607 3296 3633 3304
rect 4467 3296 4633 3304
rect 816 3276 913 3284
rect 1007 3276 1813 3284
rect 1827 3276 1953 3284
rect 1967 3276 2033 3284
rect 2287 3276 2353 3284
rect 3107 3276 3213 3284
rect 3907 3276 3913 3284
rect 3927 3276 3953 3284
rect 3987 3276 4013 3284
rect 4447 3276 4513 3284
rect 4636 3276 4673 3284
rect 127 3256 364 3264
rect 96 3227 104 3253
rect 156 3236 173 3244
rect 156 3224 164 3236
rect 356 3227 364 3256
rect 447 3256 473 3264
rect 487 3256 593 3264
rect 667 3256 813 3264
rect 856 3256 873 3264
rect 387 3236 413 3244
rect 856 3227 864 3256
rect 896 3256 953 3264
rect 896 3244 904 3256
rect 967 3256 1053 3264
rect 1067 3256 1173 3264
rect 1267 3256 1273 3264
rect 1287 3256 1364 3264
rect 1356 3247 1364 3256
rect 1507 3256 1513 3264
rect 1527 3256 1593 3264
rect 1707 3256 1824 3264
rect 887 3236 904 3244
rect 947 3236 993 3244
rect 1056 3236 1073 3244
rect 116 3216 164 3224
rect 27 3196 93 3204
rect 116 3184 124 3216
rect 187 3216 213 3224
rect 447 3216 473 3224
rect 607 3216 733 3224
rect 1056 3224 1064 3236
rect 1287 3236 1313 3244
rect 907 3216 1064 3224
rect 1087 3216 1113 3224
rect 1396 3224 1404 3253
rect 1567 3236 1613 3244
rect 1127 3216 1404 3224
rect 1447 3216 1533 3224
rect 1636 3224 1644 3253
rect 1636 3216 1693 3224
rect 1727 3216 1793 3224
rect 147 3196 233 3204
rect 247 3196 353 3204
rect 367 3196 553 3204
rect 747 3196 793 3204
rect 827 3196 833 3204
rect 847 3196 1173 3204
rect 1347 3196 1453 3204
rect 1567 3196 1713 3204
rect 1816 3204 1824 3256
rect 1907 3256 1973 3264
rect 1836 3244 1844 3253
rect 1916 3244 1924 3256
rect 2127 3256 2264 3264
rect 1836 3236 1904 3244
rect 1916 3236 2044 3244
rect 1896 3227 1904 3236
rect 2036 3227 2044 3236
rect 2076 3227 2084 3253
rect 2256 3247 2264 3256
rect 2307 3256 2404 3264
rect 2116 3236 2133 3244
rect 2116 3227 2124 3236
rect 2167 3236 2204 3244
rect 2196 3227 2204 3236
rect 1847 3216 1873 3224
rect 1816 3196 1833 3204
rect 1936 3204 1944 3213
rect 1887 3196 1944 3204
rect 2216 3204 2224 3233
rect 2247 3216 2273 3224
rect 2336 3207 2344 3233
rect 2396 3227 2404 3256
rect 3376 3256 3433 3264
rect 2967 3236 3013 3244
rect 3067 3236 3093 3244
rect 3136 3227 3144 3253
rect 3167 3236 3293 3244
rect 3307 3236 3353 3244
rect 3376 3227 3384 3256
rect 3547 3256 3613 3264
rect 3887 3256 4033 3264
rect 4156 3256 4284 3264
rect 3696 3244 3704 3253
rect 3607 3236 3704 3244
rect 3956 3236 4013 3244
rect 3956 3227 3964 3236
rect 4156 3244 4164 3256
rect 4076 3236 4164 3244
rect 2787 3216 2833 3224
rect 2847 3216 2973 3224
rect 3047 3216 3113 3224
rect 3247 3216 3313 3224
rect 3467 3216 3753 3224
rect 4076 3224 4084 3236
rect 4007 3216 4084 3224
rect 4176 3224 4184 3233
rect 4107 3216 4184 3224
rect 4207 3216 4233 3224
rect 2087 3196 2224 3204
rect 2456 3187 2464 3213
rect 4256 3207 4264 3233
rect 4276 3227 4284 3256
rect 4296 3256 4313 3264
rect 2567 3196 2853 3204
rect 3047 3196 3093 3204
rect 3187 3196 3273 3204
rect 3407 3196 3473 3204
rect 4027 3196 4113 3204
rect 4296 3204 4304 3256
rect 4416 3264 4424 3273
rect 4347 3256 4404 3264
rect 4416 3256 4473 3264
rect 4287 3196 4304 3204
rect 4376 3204 4384 3233
rect 4396 3224 4404 3256
rect 4427 3236 4493 3244
rect 4396 3216 4413 3224
rect 4347 3196 4384 3204
rect 116 3176 133 3184
rect 167 3176 313 3184
rect 347 3176 373 3184
rect 467 3176 593 3184
rect 667 3176 773 3184
rect 887 3176 1493 3184
rect 1527 3176 1993 3184
rect 2727 3176 3073 3184
rect 3987 3176 4173 3184
rect 4187 3176 4353 3184
rect 4367 3176 4433 3184
rect 4636 3184 4644 3276
rect 4656 3207 4664 3253
rect 4687 3236 4733 3244
rect 4707 3216 4733 3224
rect 4636 3176 4733 3184
rect 107 3156 393 3164
rect 467 3156 573 3164
rect 627 3156 653 3164
rect 767 3156 873 3164
rect 947 3156 973 3164
rect 1147 3156 1213 3164
rect 1247 3156 1413 3164
rect 1487 3156 1613 3164
rect 1707 3156 1773 3164
rect 1807 3156 2664 3164
rect 147 3136 293 3144
rect 647 3136 673 3144
rect 1127 3136 1393 3144
rect 1747 3136 1813 3144
rect 1927 3136 1973 3144
rect 2387 3136 2633 3144
rect 2656 3144 2664 3156
rect 2687 3156 2773 3164
rect 2907 3156 3333 3164
rect 3356 3156 3813 3164
rect 3356 3144 3364 3156
rect 3847 3156 4013 3164
rect 4067 3156 4213 3164
rect 4267 3156 4393 3164
rect 2656 3136 3364 3144
rect 3587 3136 3633 3144
rect 3927 3136 3993 3144
rect 4007 3136 4253 3144
rect 4307 3136 4373 3144
rect 247 3116 273 3124
rect 287 3116 433 3124
rect 927 3116 1213 3124
rect 1747 3116 1953 3124
rect 2167 3116 2513 3124
rect 2987 3116 3253 3124
rect 3867 3116 3993 3124
rect 4027 3116 4073 3124
rect 4247 3116 4293 3124
rect 4367 3116 4393 3124
rect 487 3096 553 3104
rect 587 3096 593 3104
rect 607 3096 784 3104
rect 76 3076 253 3084
rect 36 3007 44 3033
rect 76 3007 84 3076
rect 527 3076 593 3084
rect 776 3084 784 3096
rect 807 3096 993 3104
rect 1016 3096 1073 3104
rect 1016 3084 1024 3096
rect 1187 3096 1324 3104
rect 776 3076 1024 3084
rect 1047 3076 1193 3084
rect 1267 3076 1293 3084
rect 1316 3084 1324 3096
rect 1507 3096 1653 3104
rect 1667 3096 1753 3104
rect 1767 3096 1853 3104
rect 1887 3096 2033 3104
rect 2047 3096 2173 3104
rect 2367 3096 2713 3104
rect 2867 3096 2873 3104
rect 2887 3096 2893 3104
rect 3407 3096 3633 3104
rect 3727 3096 4113 3104
rect 4667 3096 4804 3104
rect 1316 3076 1473 3084
rect 1527 3076 1713 3084
rect 1727 3076 2093 3084
rect 2107 3076 2133 3084
rect 2287 3076 2453 3084
rect 2867 3076 3113 3084
rect 3167 3076 3373 3084
rect 3507 3076 3713 3084
rect 3787 3076 3924 3084
rect 96 3056 153 3064
rect 96 3027 104 3056
rect 356 3056 533 3064
rect -24 2964 -16 3004
rect 116 3004 124 3033
rect 276 3016 293 3024
rect 116 2996 213 3004
rect 67 2976 93 2984
rect 276 2984 284 3016
rect 356 3004 364 3056
rect 847 3056 1013 3064
rect 1187 3056 1784 3064
rect 387 3036 513 3044
rect 607 3036 724 3044
rect 547 3016 593 3024
rect 307 2996 364 3004
rect 387 2996 573 3004
rect 587 2996 673 3004
rect 276 2976 473 2984
rect 696 2984 704 3013
rect 716 3007 724 3036
rect 767 3036 833 3044
rect 1156 3044 1164 3053
rect 1156 3036 1224 3044
rect 856 3024 864 3033
rect 816 3016 864 3024
rect 976 3024 984 3033
rect 976 3016 1173 3024
rect 816 3007 824 3016
rect 947 2996 993 3004
rect 1216 3004 1224 3036
rect 1536 3036 1573 3044
rect 1276 3024 1284 3033
rect 1247 3016 1513 3024
rect 1216 2996 1253 3004
rect 1287 2996 1413 3004
rect 1427 2996 1473 3004
rect 1536 3004 1544 3036
rect 1627 3036 1753 3044
rect 1776 3027 1784 3056
rect 2127 3056 2384 3064
rect 1796 3036 1893 3044
rect 1567 3016 1704 3024
rect 1696 3007 1704 3016
rect 1796 3007 1804 3036
rect 1936 3024 1944 3053
rect 2147 3036 2193 3044
rect 2247 3036 2293 3044
rect 2336 3036 2353 3044
rect 1887 3016 1944 3024
rect 2067 3016 2073 3024
rect 2087 3016 2113 3024
rect 2167 3016 2213 3024
rect 1536 2996 1553 3004
rect 687 2976 704 2984
rect 787 2976 893 2984
rect 907 2976 1233 2984
rect 1407 2976 1453 2984
rect 1547 2976 1573 2984
rect 1816 2984 1824 3013
rect 1847 2996 1973 3004
rect 2087 2996 2293 3004
rect 1667 2976 1824 2984
rect 2316 2984 2324 3013
rect 2336 3007 2344 3036
rect 2376 3027 2384 3056
rect 2627 3056 2753 3064
rect 2767 3056 2793 3064
rect 3067 3056 3093 3064
rect 3596 3056 3673 3064
rect 2436 3044 2444 3053
rect 2396 3036 2444 3044
rect 2396 3007 2404 3036
rect 2527 3036 2653 3044
rect 2667 3036 2673 3044
rect 3087 3036 3193 3044
rect 2427 3016 2453 3024
rect 2487 3016 2533 3024
rect 2696 3004 2704 3033
rect 3036 3024 3044 3033
rect 3176 3027 3184 3036
rect 3036 3016 3153 3024
rect 3216 3024 3224 3053
rect 3367 3036 3433 3044
rect 3196 3016 3224 3024
rect 2547 2996 2704 3004
rect 2316 2976 2453 2984
rect 2716 2984 2724 3013
rect 2747 2996 2833 3004
rect 3007 2996 3033 3004
rect 3196 3004 3204 3016
rect 3507 3016 3533 3024
rect 3147 2996 3204 3004
rect 3307 2996 3393 3004
rect 2607 2976 2724 2984
rect 2987 2976 3053 2984
rect 3067 2976 3253 2984
rect 3596 2984 3604 3056
rect 3916 3064 3924 3076
rect 3987 3076 4013 3084
rect 4047 3076 4133 3084
rect 4147 3076 4313 3084
rect 4376 3076 4413 3084
rect 3916 3056 4093 3064
rect 4107 3056 4193 3064
rect 4207 3056 4233 3064
rect 4247 3056 4333 3064
rect 3647 3036 3673 3044
rect 3727 3036 3753 3044
rect 3896 3044 3904 3053
rect 3867 3036 3884 3044
rect 3896 3036 3944 3044
rect 3627 3016 3773 3024
rect 3796 3024 3804 3033
rect 3787 3016 3804 3024
rect 3827 3016 3853 3024
rect 3876 3024 3884 3036
rect 3876 3016 3893 3024
rect 3936 3024 3944 3036
rect 3967 3036 3984 3044
rect 3936 3016 3964 3024
rect 3667 2996 3713 3004
rect 3596 2976 3713 2984
rect 3956 2984 3964 3016
rect 3976 3007 3984 3036
rect 4087 3036 4144 3044
rect 4007 3016 4024 3024
rect 4016 3004 4024 3016
rect 4067 3016 4113 3024
rect 4136 3007 4144 3036
rect 4256 3036 4293 3044
rect 4176 3007 4184 3033
rect 4256 3024 4264 3036
rect 4316 3036 4353 3044
rect 4247 3016 4264 3024
rect 4276 3016 4293 3024
rect 4016 2996 4113 3004
rect 4276 2987 4284 3016
rect 4316 3004 4324 3036
rect 4376 3044 4384 3076
rect 4487 3076 4493 3084
rect 4507 3076 4633 3084
rect 4667 3076 4773 3084
rect 4407 3056 4544 3064
rect 4536 3047 4544 3056
rect 4687 3056 4733 3064
rect 4796 3064 4804 3096
rect 4787 3056 4804 3064
rect 4376 3036 4404 3044
rect 4396 3024 4404 3036
rect 4427 3036 4444 3044
rect 4396 3016 4413 3024
rect 4436 3024 4444 3036
rect 4627 3036 4673 3044
rect 4436 3016 4613 3024
rect 4707 3016 4733 3024
rect 4296 2996 4324 3004
rect 4296 2987 4304 2996
rect 4367 2996 4593 3004
rect 4607 2996 4653 3004
rect 4667 2996 4673 3004
rect 3956 2976 4093 2984
rect 4567 2976 4693 2984
rect -24 2956 373 2964
rect 447 2956 693 2964
rect 727 2956 873 2964
rect 1027 2956 1053 2964
rect 1307 2956 1593 2964
rect 1627 2956 2013 2964
rect 3387 2956 3813 2964
rect 4167 2956 4413 2964
rect 27 2936 173 2944
rect 507 2936 613 2944
rect 627 2936 753 2944
rect 967 2936 1093 2944
rect 1107 2936 1793 2944
rect 3107 2936 3433 2944
rect 4247 2936 4313 2944
rect 67 2916 313 2924
rect 567 2916 1453 2924
rect 1507 2916 1693 2924
rect 3747 2916 3773 2924
rect 4287 2916 4613 2924
rect 4627 2916 4773 2924
rect 267 2896 573 2904
rect 667 2896 873 2904
rect 896 2896 1693 2904
rect 896 2884 904 2896
rect 367 2876 904 2884
rect 1127 2876 1173 2884
rect 1367 2876 1673 2884
rect 1767 2876 3093 2884
rect 3647 2876 3833 2884
rect 3847 2876 4433 2884
rect 207 2856 1553 2864
rect 1567 2856 2773 2864
rect 2787 2856 2993 2864
rect 3687 2856 4273 2864
rect 4287 2856 4473 2864
rect 87 2836 553 2844
rect 627 2836 733 2844
rect 867 2836 893 2844
rect 907 2836 1573 2844
rect 1587 2836 1913 2844
rect 2267 2836 2953 2844
rect 3827 2836 4253 2844
rect 247 2816 273 2824
rect 567 2816 624 2824
rect 347 2796 444 2804
rect 27 2776 133 2784
rect 307 2776 353 2784
rect 387 2776 424 2784
rect -24 2684 -16 2764
rect 36 2727 44 2753
rect 56 2744 64 2753
rect 56 2736 113 2744
rect 156 2744 164 2773
rect 156 2736 173 2744
rect 196 2727 204 2753
rect 216 2724 224 2773
rect 247 2756 393 2764
rect 416 2747 424 2776
rect 436 2764 444 2796
rect 616 2804 624 2816
rect 687 2816 833 2824
rect 1067 2816 1133 2824
rect 1327 2816 1613 2824
rect 1707 2816 2493 2824
rect 3787 2816 3933 2824
rect 4047 2816 4133 2824
rect 616 2796 664 2804
rect 436 2756 493 2764
rect 267 2736 273 2744
rect 287 2736 373 2744
rect 447 2736 493 2744
rect 536 2744 544 2793
rect 576 2747 584 2773
rect 656 2764 664 2796
rect 767 2796 1193 2804
rect 1207 2796 1373 2804
rect 1387 2796 1753 2804
rect 1787 2796 1893 2804
rect 2027 2796 2053 2804
rect 2247 2796 2473 2804
rect 2507 2796 2633 2804
rect 2827 2796 3093 2804
rect 3107 2796 3853 2804
rect 4567 2796 4613 2804
rect 4627 2796 4673 2804
rect 636 2756 664 2764
rect 536 2736 553 2744
rect 636 2744 644 2756
rect 627 2736 644 2744
rect 716 2744 724 2793
rect 827 2776 953 2784
rect 1107 2776 1193 2784
rect 1267 2776 1404 2784
rect 847 2756 1004 2764
rect 687 2736 724 2744
rect 747 2736 764 2744
rect 216 2716 293 2724
rect 367 2716 533 2724
rect 756 2724 764 2736
rect 827 2736 853 2744
rect 907 2736 913 2744
rect 927 2736 973 2744
rect 996 2744 1004 2756
rect 1027 2756 1353 2764
rect 996 2736 1053 2744
rect 1087 2736 1153 2744
rect 1187 2736 1373 2744
rect 756 2716 804 2724
rect 27 2696 53 2704
rect 67 2696 213 2704
rect 347 2696 613 2704
rect 667 2696 773 2704
rect 796 2704 804 2716
rect 1027 2716 1293 2724
rect 1396 2724 1404 2776
rect 1987 2776 2213 2784
rect 2367 2776 2433 2784
rect 2487 2776 2553 2784
rect 2567 2776 2593 2784
rect 2867 2776 2913 2784
rect 3496 2776 3533 2784
rect 1636 2764 1644 2773
rect 1467 2756 1813 2764
rect 1836 2747 1844 2773
rect 1867 2756 1893 2764
rect 1947 2756 2153 2764
rect 2216 2756 2273 2764
rect 1867 2736 1993 2744
rect 2216 2744 2224 2756
rect 2347 2756 2373 2764
rect 2556 2756 2633 2764
rect 2147 2736 2224 2744
rect 2416 2744 2424 2753
rect 2556 2747 2564 2756
rect 2787 2756 2833 2764
rect 2416 2736 2433 2744
rect 2527 2736 2553 2744
rect 2736 2744 2744 2753
rect 3496 2747 3504 2776
rect 3567 2776 3593 2784
rect 3607 2776 3653 2784
rect 3807 2776 3893 2784
rect 3956 2776 4144 2784
rect 2587 2736 2744 2744
rect 2767 2736 2973 2744
rect 3607 2736 3653 2744
rect 3956 2744 3964 2776
rect 4136 2767 4144 2776
rect 4196 2776 4213 2784
rect 3987 2756 4024 2764
rect 3887 2736 3964 2744
rect 4016 2744 4024 2756
rect 4196 2764 4204 2776
rect 4507 2776 4633 2784
rect 4176 2756 4204 2764
rect 4016 2736 4044 2744
rect 1316 2716 1404 2724
rect 1756 2724 1764 2733
rect 1756 2716 1893 2724
rect 796 2696 1033 2704
rect 1047 2696 1113 2704
rect 1127 2696 1213 2704
rect 1316 2704 1324 2716
rect 1907 2716 2093 2724
rect 2207 2716 2253 2724
rect 2267 2716 2313 2724
rect 2667 2716 2713 2724
rect 2887 2716 3013 2724
rect 3027 2716 3253 2724
rect 3427 2716 3433 2724
rect 3447 2716 3833 2724
rect 3987 2716 4013 2724
rect 4036 2724 4044 2736
rect 4176 2744 4184 2756
rect 4636 2747 4644 2773
rect 4067 2736 4184 2744
rect 4387 2736 4573 2744
rect 4687 2736 4753 2744
rect 4036 2716 4053 2724
rect 4127 2716 4173 2724
rect 4207 2716 4233 2724
rect 4287 2716 4413 2724
rect 4447 2716 4533 2724
rect 4607 2716 4653 2724
rect 1267 2696 1324 2704
rect 1647 2696 1853 2704
rect 1967 2696 2053 2704
rect 2287 2696 2453 2704
rect 2467 2696 2533 2704
rect 2727 2696 2793 2704
rect 3127 2696 3213 2704
rect 3507 2696 3733 2704
rect 3747 2696 3853 2704
rect 3867 2696 3893 2704
rect 3947 2696 3993 2704
rect 4087 2696 4113 2704
rect 4247 2696 4313 2704
rect 4567 2696 4693 2704
rect -24 2676 1133 2684
rect 1147 2676 1473 2684
rect 1496 2676 1693 2684
rect 67 2656 93 2664
rect 107 2656 313 2664
rect 427 2656 813 2664
rect 847 2656 973 2664
rect 1107 2656 1313 2664
rect 1496 2664 1504 2676
rect 1787 2676 1913 2684
rect 2047 2676 2093 2684
rect 2127 2676 2293 2684
rect 2307 2676 2633 2684
rect 3047 2676 3213 2684
rect 3227 2676 3453 2684
rect 4167 2676 4513 2684
rect 1347 2656 1504 2664
rect 1667 2656 1833 2664
rect 2287 2656 2513 2664
rect 3167 2656 3533 2664
rect 3807 2656 4133 2664
rect 807 2636 933 2644
rect 1007 2636 1133 2644
rect 1167 2636 1233 2644
rect 1687 2636 2073 2644
rect 2207 2636 2293 2644
rect 2307 2636 2393 2644
rect 3007 2636 3453 2644
rect 3487 2636 3613 2644
rect 4007 2636 4213 2644
rect 4227 2636 4393 2644
rect 107 2616 173 2624
rect 187 2616 353 2624
rect 447 2616 613 2624
rect 807 2616 853 2624
rect 867 2616 1033 2624
rect 1307 2616 1653 2624
rect 3307 2616 3533 2624
rect 3787 2616 3973 2624
rect 4067 2616 4153 2624
rect 167 2596 253 2604
rect 267 2596 553 2604
rect 47 2576 133 2584
rect 27 2556 73 2564
rect 87 2556 144 2564
rect 67 2536 113 2544
rect 136 2544 144 2556
rect 256 2556 393 2564
rect 256 2547 264 2556
rect 416 2547 424 2596
rect 567 2596 593 2604
rect 967 2596 1093 2604
rect 1187 2596 1233 2604
rect 1347 2596 1493 2604
rect 1507 2596 1593 2604
rect 1607 2596 1793 2604
rect 2387 2596 2693 2604
rect 3247 2596 3473 2604
rect 3687 2596 3813 2604
rect 3827 2596 3913 2604
rect 4027 2596 4093 2604
rect 527 2576 613 2584
rect 927 2576 953 2584
rect 987 2576 1193 2584
rect 1247 2576 1373 2584
rect 1467 2576 1493 2584
rect 1987 2576 2073 2584
rect 2087 2576 2133 2584
rect 2267 2576 2333 2584
rect 2347 2576 2464 2584
rect 456 2564 464 2573
rect 456 2556 564 2564
rect 136 2536 153 2544
rect 167 2536 233 2544
rect 447 2536 533 2544
rect 327 2516 353 2524
rect 367 2516 373 2524
rect 467 2516 533 2524
rect 556 2524 564 2556
rect 556 2516 613 2524
rect 716 2524 724 2573
rect 847 2556 864 2564
rect 707 2516 724 2524
rect 767 2516 833 2524
rect 856 2524 864 2556
rect 907 2556 964 2564
rect 887 2536 904 2544
rect 856 2516 873 2524
rect 27 2496 573 2504
rect 896 2504 904 2536
rect 956 2527 964 2556
rect 1007 2556 1013 2564
rect 1067 2556 1273 2564
rect 996 2527 1004 2553
rect 1167 2536 1184 2544
rect 1087 2516 1153 2524
rect 1176 2524 1184 2536
rect 1176 2516 1193 2524
rect 896 2496 933 2504
rect 987 2496 1133 2504
rect 1356 2504 1364 2553
rect 1436 2547 1444 2573
rect 1707 2556 1733 2564
rect 2456 2564 2464 2576
rect 2487 2576 2833 2584
rect 2847 2576 2853 2584
rect 2907 2576 3033 2584
rect 3047 2576 3333 2584
rect 3967 2576 3984 2584
rect 2456 2556 2493 2564
rect 2687 2556 2733 2564
rect 2747 2556 2793 2564
rect 2927 2556 3073 2564
rect 3087 2556 3193 2564
rect 1476 2524 1484 2553
rect 1547 2536 1633 2544
rect 1476 2516 1513 2524
rect 1567 2516 1593 2524
rect 1607 2516 1653 2524
rect 1667 2516 1813 2524
rect 1287 2496 1364 2504
rect 1407 2496 1413 2504
rect 1427 2496 1593 2504
rect 1827 2496 1893 2504
rect 1936 2504 1944 2553
rect 2027 2536 2093 2544
rect 2116 2544 2124 2553
rect 2107 2536 2124 2544
rect 2187 2536 2193 2544
rect 2207 2536 2213 2544
rect 2327 2536 2373 2544
rect 2007 2516 2053 2524
rect 2396 2524 2404 2553
rect 2427 2536 2693 2544
rect 2787 2536 2924 2544
rect 2916 2527 2924 2536
rect 2947 2536 3093 2544
rect 3147 2536 3293 2544
rect 3356 2544 3364 2573
rect 3487 2556 3593 2564
rect 3707 2556 3873 2564
rect 3356 2536 3393 2544
rect 3787 2536 3893 2544
rect 3956 2544 3964 2553
rect 3976 2547 3984 2576
rect 4087 2576 4473 2584
rect 4007 2556 4033 2564
rect 4327 2556 4513 2564
rect 4547 2556 4593 2564
rect 3947 2536 3964 2544
rect 4207 2536 4213 2544
rect 4227 2536 4333 2544
rect 4447 2536 4584 2544
rect 4576 2527 4584 2536
rect 4616 2527 4624 2553
rect 2347 2516 2404 2524
rect 2587 2516 2793 2524
rect 2807 2516 2853 2524
rect 3327 2516 3393 2524
rect 3447 2516 3513 2524
rect 3527 2516 4053 2524
rect 4267 2516 4313 2524
rect 4447 2516 4553 2524
rect 4647 2516 4693 2524
rect 1936 2496 2033 2504
rect 2567 2496 2573 2504
rect 2587 2496 2653 2504
rect 2727 2496 2813 2504
rect 2887 2496 2953 2504
rect 3287 2496 3553 2504
rect 3567 2496 3573 2504
rect 3827 2496 4033 2504
rect 4047 2496 4093 2504
rect 4467 2496 4653 2504
rect 487 2476 593 2484
rect 727 2476 813 2484
rect 827 2476 833 2484
rect 967 2476 1013 2484
rect 1367 2476 1413 2484
rect 1427 2476 1673 2484
rect 1807 2476 1853 2484
rect 1967 2476 2033 2484
rect 3867 2476 3933 2484
rect 3967 2476 4233 2484
rect 4507 2476 4613 2484
rect 4627 2476 4693 2484
rect 347 2456 773 2464
rect 927 2456 1113 2464
rect 1827 2456 2093 2464
rect 3267 2456 4073 2464
rect 987 2436 1073 2444
rect 4067 2436 4113 2444
rect 427 2416 493 2424
rect 587 2416 1433 2424
rect 1787 2416 1933 2424
rect 1947 2416 2153 2424
rect 2927 2416 2973 2424
rect 47 2396 213 2404
rect 767 2396 813 2404
rect 827 2396 873 2404
rect 1047 2396 1253 2404
rect 3787 2396 4013 2404
rect 687 2376 993 2384
rect 1007 2376 1153 2384
rect 1507 2376 1633 2384
rect 3827 2376 3993 2384
rect 147 2356 273 2364
rect 327 2356 453 2364
rect 767 2356 1473 2364
rect 2267 2356 2633 2364
rect 3107 2356 3533 2364
rect 3587 2356 3673 2364
rect 3707 2356 3873 2364
rect 76 2336 413 2344
rect 16 2224 24 2313
rect 36 2267 44 2313
rect 76 2284 84 2336
rect 96 2287 104 2313
rect 207 2296 293 2304
rect 316 2287 324 2313
rect 67 2276 84 2284
rect 107 2276 164 2284
rect 87 2256 133 2264
rect 156 2264 164 2276
rect 187 2276 233 2284
rect 287 2276 313 2284
rect 336 2284 344 2336
rect 967 2336 1193 2344
rect 1327 2336 1353 2344
rect 1487 2336 1573 2344
rect 2527 2336 2673 2344
rect 3956 2336 4133 2344
rect 527 2316 633 2324
rect 1127 2316 1133 2324
rect 1147 2316 1313 2324
rect 2287 2316 2613 2324
rect 356 2304 364 2313
rect 356 2296 384 2304
rect 336 2276 353 2284
rect 376 2267 384 2296
rect 667 2296 733 2304
rect 856 2296 913 2304
rect 156 2256 333 2264
rect 436 2264 444 2273
rect 436 2256 464 2264
rect 207 2236 213 2244
rect 227 2236 293 2244
rect 347 2236 433 2244
rect 456 2244 464 2256
rect 536 2264 544 2273
rect 487 2256 544 2264
rect 567 2256 593 2264
rect 456 2236 473 2244
rect 676 2227 684 2273
rect 696 2264 704 2273
rect 856 2267 864 2296
rect 1007 2296 1093 2304
rect 1107 2296 1253 2304
rect 1987 2296 2073 2304
rect 2367 2296 2393 2304
rect 2536 2304 2544 2316
rect 3307 2316 3633 2324
rect 3667 2316 3713 2324
rect 2527 2296 2544 2304
rect 2567 2296 2613 2304
rect 3007 2296 3153 2304
rect 3567 2296 3773 2304
rect 956 2267 964 2293
rect 1047 2276 1173 2284
rect 1567 2276 1613 2284
rect 1927 2276 1973 2284
rect 2027 2276 2213 2284
rect 2267 2276 2324 2284
rect 696 2256 793 2264
rect 927 2256 953 2264
rect 1027 2256 1053 2264
rect 1067 2256 1073 2264
rect 1216 2264 1224 2273
rect 2316 2267 2324 2276
rect 2387 2276 2433 2284
rect 2487 2276 2533 2284
rect 2867 2276 3084 2284
rect 1187 2256 1224 2264
rect 1247 2256 1384 2264
rect 847 2236 953 2244
rect 987 2236 1093 2244
rect 1207 2236 1333 2244
rect 1376 2244 1384 2256
rect 1427 2256 1453 2264
rect 1587 2256 1653 2264
rect 1807 2256 2244 2264
rect 1376 2236 1573 2244
rect 1847 2236 1913 2244
rect 2236 2244 2244 2256
rect 2267 2256 2293 2264
rect 2376 2247 2384 2273
rect 3076 2267 3084 2276
rect 3176 2276 3493 2284
rect 3176 2267 3184 2276
rect 3596 2276 3613 2284
rect 3596 2267 3604 2276
rect 3667 2276 3684 2284
rect 3676 2267 3684 2276
rect 3727 2276 3784 2284
rect 3776 2267 3784 2276
rect 3816 2267 3824 2293
rect 2427 2256 2573 2264
rect 2807 2256 2933 2264
rect 2987 2256 3053 2264
rect 3207 2256 3233 2264
rect 3247 2256 3253 2264
rect 3387 2256 3513 2264
rect 3647 2256 3673 2264
rect 3916 2264 3924 2273
rect 3936 2267 3944 2293
rect 3956 2287 3964 2336
rect 4587 2336 4773 2344
rect 3987 2316 4084 2324
rect 4016 2296 4053 2304
rect 4016 2267 4024 2296
rect 3836 2256 3924 2264
rect 2236 2236 2264 2244
rect 2256 2227 2264 2236
rect 2287 2236 2353 2244
rect 2547 2236 2613 2244
rect 2947 2236 3333 2244
rect 3347 2236 3493 2244
rect 3607 2236 3653 2244
rect 3836 2244 3844 2256
rect 3947 2256 4004 2264
rect 3996 2247 4004 2256
rect 3727 2236 3844 2244
rect 3867 2236 3973 2244
rect 4036 2244 4044 2273
rect 4016 2236 4044 2244
rect 4016 2227 4024 2236
rect 16 2216 213 2224
rect 247 2216 273 2224
rect 407 2216 513 2224
rect 527 2216 573 2224
rect 847 2216 933 2224
rect 987 2216 1133 2224
rect 1167 2216 1253 2224
rect 1547 2216 1673 2224
rect 1887 2216 1953 2224
rect 1967 2216 2113 2224
rect 2176 2216 2193 2224
rect 167 2196 353 2204
rect 367 2196 553 2204
rect 567 2196 653 2204
rect 827 2196 913 2204
rect 1387 2196 1713 2204
rect 1827 2196 1933 2204
rect 2176 2187 2184 2216
rect 2667 2216 3213 2224
rect 3367 2216 3513 2224
rect 4076 2224 4084 2316
rect 4587 2316 4693 2324
rect 4347 2296 4533 2304
rect 4547 2296 4653 2304
rect 4627 2276 4673 2284
rect 4227 2256 4413 2264
rect 4467 2256 4593 2264
rect 4687 2256 4733 2264
rect 4167 2236 4233 2244
rect 4047 2216 4084 2224
rect 2467 2196 2693 2204
rect 2707 2196 2953 2204
rect 3127 2196 3293 2204
rect 3607 2196 3753 2204
rect 3767 2196 3833 2204
rect 27 2176 313 2184
rect 587 2176 713 2184
rect 1647 2176 1693 2184
rect 1787 2176 1993 2184
rect 2907 2176 2973 2184
rect 2987 2176 3013 2184
rect 3027 2176 3133 2184
rect 3147 2176 3173 2184
rect 3587 2176 4553 2184
rect 287 2156 533 2164
rect 547 2156 893 2164
rect 1707 2156 1813 2164
rect 1847 2156 1873 2164
rect 1947 2156 2233 2164
rect 2547 2156 2593 2164
rect 2607 2156 2673 2164
rect 2927 2156 3253 2164
rect 4547 2156 4593 2164
rect 187 2136 753 2144
rect 1327 2136 1753 2144
rect 1767 2136 2053 2144
rect 2167 2136 2293 2144
rect 2667 2136 3273 2144
rect 3687 2136 3793 2144
rect 3827 2136 3933 2144
rect 4307 2136 4373 2144
rect 4427 2136 4533 2144
rect 4547 2136 4633 2144
rect 467 2116 573 2124
rect 647 2116 713 2124
rect 736 2116 793 2124
rect 36 2096 53 2104
rect 36 2044 44 2096
rect 87 2096 324 2104
rect 67 2076 133 2084
rect 156 2076 173 2084
rect 156 2064 164 2076
rect 267 2076 304 2084
rect 96 2056 164 2064
rect 96 2047 104 2056
rect 36 2036 73 2044
rect 216 2044 224 2073
rect 187 2036 224 2044
rect 236 2027 244 2073
rect 296 2067 304 2076
rect 316 2067 324 2096
rect 367 2096 404 2104
rect 367 2076 384 2084
rect 276 2044 284 2053
rect 276 2036 333 2044
rect 376 2044 384 2076
rect 396 2067 404 2096
rect 416 2096 473 2104
rect 416 2067 424 2096
rect 736 2104 744 2116
rect 947 2116 1033 2124
rect 1667 2116 1893 2124
rect 1927 2116 1973 2124
rect 2067 2116 2213 2124
rect 3007 2116 3033 2124
rect 3207 2116 3244 2124
rect 496 2096 744 2104
rect 496 2084 504 2096
rect 807 2096 884 2104
rect 436 2076 504 2084
rect 436 2067 444 2076
rect 776 2084 784 2093
rect 756 2076 784 2084
rect 796 2076 813 2084
rect 536 2056 593 2064
rect 376 2036 393 2044
rect 447 2036 513 2044
rect 256 2004 264 2033
rect 536 2024 544 2056
rect 656 2064 664 2073
rect 656 2056 693 2064
rect 636 2044 644 2053
rect 756 2047 764 2076
rect 567 2036 713 2044
rect 796 2044 804 2076
rect 876 2084 884 2096
rect 907 2096 1013 2104
rect 1127 2096 1213 2104
rect 1236 2096 1413 2104
rect 876 2076 933 2084
rect 1007 2076 1064 2084
rect 827 2056 913 2064
rect 796 2036 873 2044
rect 956 2044 964 2073
rect 1027 2056 1044 2064
rect 936 2036 964 2044
rect 536 2016 564 2024
rect 27 1996 264 2004
rect 276 1996 513 2004
rect 276 1984 284 1996
rect 556 2004 564 2016
rect 647 2016 793 2024
rect 916 2024 924 2033
rect 936 2027 944 2036
rect 907 2016 924 2024
rect 1016 2024 1024 2033
rect 1036 2027 1044 2056
rect 1056 2027 1064 2076
rect 1116 2076 1153 2084
rect 1096 2027 1104 2053
rect 1007 2016 1024 2024
rect 1116 2024 1124 2076
rect 1147 2056 1193 2064
rect 1236 2064 1244 2096
rect 1867 2096 1933 2104
rect 2287 2096 2393 2104
rect 2407 2096 2573 2104
rect 3067 2096 3213 2104
rect 1267 2076 1293 2084
rect 1347 2076 1373 2084
rect 1567 2076 1693 2084
rect 1736 2067 1744 2093
rect 1756 2067 1764 2093
rect 1956 2084 1964 2093
rect 1936 2076 1964 2084
rect 1227 2056 1244 2064
rect 1287 2056 1313 2064
rect 1507 2056 1633 2064
rect 1687 2056 1713 2064
rect 1167 2036 1433 2044
rect 1447 2036 1533 2044
rect 1116 2016 1293 2024
rect 1407 2016 1733 2024
rect 1747 2016 1893 2024
rect 1916 2024 1924 2073
rect 1936 2047 1944 2076
rect 2047 2076 2113 2084
rect 2567 2076 2673 2084
rect 2927 2076 3093 2084
rect 3156 2076 3173 2084
rect 3156 2067 3164 2076
rect 3236 2084 3244 2116
rect 3547 2116 4313 2124
rect 4327 2116 4473 2124
rect 3627 2096 3813 2104
rect 3847 2096 4053 2104
rect 4067 2096 4193 2104
rect 4367 2096 4413 2104
rect 3196 2076 3244 2084
rect 1967 2056 2093 2064
rect 2347 2056 2413 2064
rect 2727 2056 2764 2064
rect 2756 2047 2764 2056
rect 2787 2056 3133 2064
rect 3196 2064 3204 2076
rect 3327 2076 3453 2084
rect 3547 2076 3573 2084
rect 3667 2076 3793 2084
rect 3887 2076 3973 2084
rect 3987 2076 4033 2084
rect 4336 2084 4344 2093
rect 4316 2076 4344 2084
rect 3176 2056 3204 2064
rect 2687 2036 2733 2044
rect 2807 2036 2913 2044
rect 3176 2044 3184 2056
rect 3267 2056 3293 2064
rect 3616 2064 3624 2073
rect 3347 2056 3624 2064
rect 4096 2064 4104 2073
rect 4316 2067 4324 2076
rect 4496 2067 4504 2093
rect 4527 2076 4553 2084
rect 3927 2056 4104 2064
rect 4347 2056 4373 2064
rect 3127 2036 3184 2044
rect 3387 2036 4333 2044
rect 1916 2016 1993 2024
rect 3447 2016 3493 2024
rect 3807 2016 3813 2024
rect 3827 2016 4053 2024
rect 556 1996 733 2004
rect 787 1996 853 2004
rect 987 1996 1073 2004
rect 1127 1996 1173 2004
rect 1527 1996 1573 2004
rect 1887 1996 2013 2004
rect 2627 1996 2693 2004
rect 2707 1996 2753 2004
rect 3147 1996 3633 2004
rect 187 1976 284 1984
rect 667 1976 893 1984
rect 907 1976 993 1984
rect 1367 1976 1653 1984
rect 1927 1976 2233 1984
rect 2387 1976 2653 1984
rect 227 1956 693 1964
rect 707 1956 853 1964
rect 2527 1956 2673 1964
rect 4007 1956 4073 1964
rect 247 1936 293 1944
rect 2087 1936 2093 1944
rect 2107 1936 2153 1944
rect 2167 1936 2393 1944
rect 2827 1936 3273 1944
rect 3627 1936 3713 1944
rect 3907 1936 4013 1944
rect 4167 1936 4193 1944
rect 247 1916 553 1924
rect 687 1916 773 1924
rect 1407 1916 1453 1924
rect 4207 1916 4233 1924
rect 327 1896 613 1904
rect 727 1896 1013 1904
rect 1727 1896 1753 1904
rect 27 1876 93 1884
rect 407 1876 833 1884
rect 847 1876 893 1884
rect 967 1876 1433 1884
rect 47 1856 213 1864
rect 307 1856 373 1864
rect 387 1856 453 1864
rect 587 1856 813 1864
rect 887 1856 953 1864
rect 1047 1856 1153 1864
rect 2207 1856 2393 1864
rect 2407 1856 2933 1864
rect 2947 1856 3153 1864
rect 3167 1856 3553 1864
rect 3667 1856 4113 1864
rect 127 1836 233 1844
rect 316 1836 413 1844
rect 56 1764 64 1833
rect 107 1816 213 1824
rect 316 1824 324 1836
rect 487 1836 713 1844
rect 867 1836 984 1844
rect 227 1816 324 1824
rect 387 1816 433 1824
rect 447 1816 573 1824
rect 587 1816 673 1824
rect 747 1816 804 1824
rect 76 1787 84 1813
rect 167 1796 184 1804
rect 176 1784 184 1796
rect 207 1796 253 1804
rect 336 1787 344 1813
rect 796 1807 804 1816
rect 827 1816 864 1824
rect 687 1796 724 1804
rect 176 1776 273 1784
rect 387 1776 453 1784
rect 507 1776 533 1784
rect 627 1776 693 1784
rect 716 1784 724 1796
rect 716 1776 733 1784
rect 56 1756 93 1764
rect 267 1756 353 1764
rect 376 1756 533 1764
rect 47 1736 173 1744
rect 376 1744 384 1756
rect 547 1756 593 1764
rect 796 1764 804 1793
rect 856 1787 864 1816
rect 827 1776 844 1784
rect 647 1756 784 1764
rect 796 1756 813 1764
rect 227 1736 384 1744
rect 427 1736 513 1744
rect 596 1736 653 1744
rect 27 1716 133 1724
rect 327 1716 393 1724
rect 596 1724 604 1736
rect 667 1736 753 1744
rect 776 1744 784 1756
rect 836 1764 844 1776
rect 867 1776 873 1784
rect 836 1756 853 1764
rect 916 1764 924 1813
rect 976 1807 984 1836
rect 996 1836 1013 1844
rect 996 1827 1004 1836
rect 1047 1836 1084 1844
rect 1076 1824 1084 1836
rect 1107 1836 1233 1844
rect 1076 1816 1093 1824
rect 1036 1787 1044 1813
rect 947 1776 1013 1784
rect 887 1756 924 1764
rect 1056 1764 1064 1813
rect 1136 1787 1144 1836
rect 1307 1836 1713 1844
rect 2167 1836 2273 1844
rect 2367 1836 2473 1844
rect 2716 1836 2733 1844
rect 1167 1816 1253 1824
rect 1276 1784 1284 1833
rect 1307 1816 1404 1824
rect 1396 1804 1404 1816
rect 1447 1816 1533 1824
rect 1627 1816 1673 1824
rect 1807 1816 1933 1824
rect 2087 1816 2193 1824
rect 2347 1816 2384 1824
rect 2376 1807 2384 1816
rect 1396 1796 1424 1804
rect 1416 1787 1424 1796
rect 1487 1796 1533 1804
rect 1567 1796 1633 1804
rect 1727 1796 1793 1804
rect 2187 1796 2253 1804
rect 2287 1796 2333 1804
rect 1276 1776 1293 1784
rect 1427 1776 1513 1784
rect 1747 1776 1813 1784
rect 1827 1776 1853 1784
rect 2147 1776 2193 1784
rect 2336 1784 2344 1793
rect 2336 1776 2493 1784
rect 2596 1784 2604 1793
rect 2547 1776 2604 1784
rect 2636 1784 2644 1793
rect 2636 1776 2693 1784
rect 1056 1756 1073 1764
rect 1087 1756 1233 1764
rect 1507 1756 1633 1764
rect 1787 1756 1833 1764
rect 2227 1756 2413 1764
rect 2507 1756 2573 1764
rect 2716 1764 2724 1836
rect 3307 1836 3333 1844
rect 3347 1836 3453 1844
rect 3467 1836 3813 1844
rect 3827 1836 4273 1844
rect 4527 1836 4553 1844
rect 2747 1816 2804 1824
rect 2796 1804 2804 1816
rect 3067 1816 3133 1824
rect 3427 1816 3513 1824
rect 3967 1816 3984 1824
rect 2796 1796 2853 1804
rect 2796 1784 2804 1796
rect 2907 1796 2953 1804
rect 3387 1796 3433 1804
rect 3867 1796 3913 1804
rect 3976 1804 3984 1816
rect 4667 1816 4733 1824
rect 3976 1796 4064 1804
rect 2787 1776 2804 1784
rect 2887 1776 2913 1784
rect 3067 1776 3073 1784
rect 3087 1776 3093 1784
rect 3336 1784 3344 1793
rect 3336 1776 3373 1784
rect 3787 1776 3813 1784
rect 3956 1784 3964 1793
rect 3887 1776 3964 1784
rect 3987 1776 4033 1784
rect 4056 1767 4064 1796
rect 4116 1796 4213 1804
rect 4116 1787 4124 1796
rect 4307 1796 4353 1804
rect 4396 1796 4453 1804
rect 2716 1756 2793 1764
rect 2827 1756 2833 1764
rect 2847 1756 3033 1764
rect 3467 1756 3493 1764
rect 3587 1756 3733 1764
rect 3767 1756 3813 1764
rect 3827 1756 4033 1764
rect 4256 1764 4264 1793
rect 4396 1784 4404 1796
rect 4347 1776 4404 1784
rect 4427 1776 4493 1784
rect 4587 1776 4673 1784
rect 4247 1756 4393 1764
rect 776 1736 913 1744
rect 967 1736 1013 1744
rect 1047 1736 1173 1744
rect 1187 1736 1273 1744
rect 1467 1736 1653 1744
rect 2367 1736 2413 1744
rect 2467 1736 2513 1744
rect 3367 1736 3633 1744
rect 3887 1736 3993 1744
rect 4087 1736 4233 1744
rect 4407 1736 4593 1744
rect 476 1716 604 1724
rect 127 1696 253 1704
rect 287 1696 453 1704
rect 476 1704 484 1716
rect 667 1716 813 1724
rect 867 1716 1253 1724
rect 1387 1716 1833 1724
rect 1847 1716 2293 1724
rect 3487 1716 3573 1724
rect 3807 1716 3953 1724
rect 4027 1716 4453 1724
rect 4467 1716 4653 1724
rect 467 1696 484 1704
rect 767 1696 933 1704
rect 1287 1696 1313 1704
rect 1327 1696 1693 1704
rect 3147 1696 3253 1704
rect 3867 1696 4073 1704
rect 4087 1696 4093 1704
rect 4227 1696 4273 1704
rect 4347 1696 4473 1704
rect 147 1676 973 1684
rect 1267 1676 1293 1684
rect 1336 1676 1613 1684
rect 367 1656 633 1664
rect 1336 1664 1344 1676
rect 2487 1676 2553 1684
rect 2787 1676 2833 1684
rect 3627 1676 3793 1684
rect 3907 1676 4293 1684
rect 4427 1676 4653 1684
rect 1147 1656 1344 1664
rect 1367 1656 1853 1664
rect 2567 1656 3333 1664
rect 3847 1656 3893 1664
rect 4067 1656 4093 1664
rect 4127 1656 4153 1664
rect 4167 1656 4273 1664
rect 4327 1656 4413 1664
rect 4447 1656 4533 1664
rect 287 1636 413 1644
rect 507 1636 573 1644
rect 587 1636 593 1644
rect 727 1636 773 1644
rect 927 1636 993 1644
rect 1127 1636 1473 1644
rect 1487 1636 1533 1644
rect 1547 1636 1573 1644
rect 1967 1636 2033 1644
rect 2167 1636 2353 1644
rect 2447 1636 2613 1644
rect 2627 1636 2673 1644
rect 2687 1636 2713 1644
rect 2767 1636 2933 1644
rect 107 1616 124 1624
rect 27 1596 93 1604
rect 116 1604 124 1616
rect 147 1616 173 1624
rect 307 1616 473 1624
rect 496 1616 533 1624
rect 116 1596 144 1604
rect 136 1587 144 1596
rect 387 1596 424 1604
rect 416 1587 424 1596
rect 496 1604 504 1616
rect 647 1616 713 1624
rect 827 1616 913 1624
rect 967 1616 1164 1624
rect 476 1596 504 1604
rect 596 1596 653 1604
rect 47 1576 113 1584
rect 167 1576 213 1584
rect 227 1576 293 1584
rect 307 1576 373 1584
rect 436 1567 444 1593
rect 476 1584 484 1596
rect 456 1576 484 1584
rect 127 1556 193 1564
rect 456 1544 464 1576
rect 596 1584 604 1596
rect 776 1596 793 1604
rect 587 1576 604 1584
rect 627 1576 693 1584
rect 776 1584 784 1596
rect 887 1596 904 1604
rect 727 1576 784 1584
rect 807 1576 813 1584
rect 847 1576 873 1584
rect 896 1584 904 1596
rect 1027 1596 1044 1604
rect 896 1576 913 1584
rect 947 1576 1013 1584
rect 796 1564 804 1573
rect 707 1556 804 1564
rect 867 1556 884 1564
rect 327 1536 464 1544
rect 616 1544 624 1553
rect 547 1536 624 1544
rect 816 1544 824 1553
rect 876 1544 884 1556
rect 907 1556 1013 1564
rect 1036 1547 1044 1596
rect 1156 1587 1164 1616
rect 1347 1616 1373 1624
rect 1547 1616 1593 1624
rect 1687 1616 1784 1624
rect 1187 1596 1193 1604
rect 1316 1604 1324 1613
rect 1207 1596 1264 1604
rect 1316 1596 1444 1604
rect 1076 1576 1113 1584
rect 1076 1564 1084 1576
rect 1196 1576 1213 1584
rect 1067 1556 1084 1564
rect 1107 1556 1153 1564
rect 1196 1564 1204 1576
rect 1256 1584 1264 1596
rect 1256 1576 1333 1584
rect 1347 1576 1413 1584
rect 1187 1556 1204 1564
rect 667 1536 864 1544
rect 876 1536 993 1544
rect 567 1516 733 1524
rect 856 1524 864 1536
rect 1216 1544 1224 1553
rect 1236 1547 1244 1573
rect 1287 1556 1333 1564
rect 1436 1564 1444 1596
rect 1627 1596 1753 1604
rect 1507 1576 1553 1584
rect 1587 1576 1673 1584
rect 1776 1584 1784 1616
rect 1756 1576 1784 1584
rect 1796 1616 1833 1624
rect 1427 1556 1444 1564
rect 1527 1556 1633 1564
rect 1207 1536 1224 1544
rect 1696 1544 1704 1573
rect 1756 1567 1764 1576
rect 1796 1567 1804 1616
rect 2027 1616 2153 1624
rect 2187 1616 2433 1624
rect 2607 1616 2733 1624
rect 1847 1596 1873 1604
rect 1816 1564 1824 1593
rect 1916 1587 1924 1613
rect 1936 1584 1944 1613
rect 2027 1596 2093 1604
rect 2207 1596 2533 1604
rect 2236 1587 2244 1596
rect 2576 1596 2633 1604
rect 2576 1587 2584 1596
rect 2707 1596 2753 1604
rect 1936 1576 1953 1584
rect 2067 1576 2113 1584
rect 2816 1584 2824 1636
rect 3147 1636 3213 1644
rect 3327 1636 3513 1644
rect 3667 1636 3744 1644
rect 2847 1616 2933 1624
rect 3007 1616 3353 1624
rect 3407 1616 3533 1624
rect 2836 1587 2844 1613
rect 2867 1596 2893 1604
rect 2927 1596 2944 1604
rect 2807 1576 2824 1584
rect 2936 1584 2944 1596
rect 2967 1596 3064 1604
rect 3056 1587 3064 1596
rect 3107 1596 3173 1604
rect 3347 1596 3384 1604
rect 2887 1576 2993 1584
rect 3067 1576 3113 1584
rect 3167 1576 3213 1584
rect 1816 1556 1833 1564
rect 1907 1556 1973 1564
rect 2007 1556 2033 1564
rect 2107 1556 2173 1564
rect 2187 1556 2333 1564
rect 2536 1564 2544 1573
rect 3236 1567 3244 1593
rect 3376 1587 3384 1596
rect 3447 1596 3473 1604
rect 3576 1567 3584 1613
rect 3736 1604 3744 1636
rect 3787 1636 4624 1644
rect 3767 1616 3864 1624
rect 3736 1596 3784 1604
rect 3776 1567 3784 1596
rect 3816 1596 3833 1604
rect 3816 1584 3824 1596
rect 3807 1576 3824 1584
rect 3856 1584 3864 1616
rect 3876 1587 3884 1636
rect 3947 1616 4073 1624
rect 3996 1607 4004 1616
rect 4267 1616 4333 1624
rect 4527 1616 4573 1624
rect 4096 1604 4104 1613
rect 4076 1596 4104 1604
rect 4176 1604 4184 1613
rect 4356 1604 4364 1613
rect 4176 1596 4244 1604
rect 3847 1576 3864 1584
rect 4076 1584 4084 1596
rect 4027 1576 4084 1584
rect 4107 1576 4213 1584
rect 4236 1584 4244 1596
rect 4336 1596 4364 1604
rect 4236 1576 4253 1584
rect 2347 1556 2553 1564
rect 2627 1556 2653 1564
rect 2787 1556 2893 1564
rect 3347 1556 3413 1564
rect 3827 1556 4313 1564
rect 4336 1564 4344 1596
rect 4387 1596 4513 1604
rect 4367 1576 4433 1584
rect 4596 1584 4604 1593
rect 4616 1587 4624 1636
rect 4647 1596 4673 1604
rect 4727 1596 4753 1604
rect 4787 1596 4804 1604
rect 4507 1576 4604 1584
rect 4727 1576 4773 1584
rect 4336 1556 4353 1564
rect 4467 1556 4473 1564
rect 4487 1556 4693 1564
rect 4796 1564 4804 1596
rect 4747 1556 4804 1564
rect 1267 1536 1704 1544
rect 1787 1536 1853 1544
rect 2127 1536 2373 1544
rect 2807 1536 2913 1544
rect 3187 1536 3193 1544
rect 3207 1536 3333 1544
rect 3487 1536 3713 1544
rect 4067 1536 4133 1544
rect 4207 1536 4253 1544
rect 856 1516 893 1524
rect 1307 1516 1613 1524
rect 3307 1516 3353 1524
rect 4387 1516 4633 1524
rect 487 1496 693 1504
rect 807 1496 913 1504
rect 1007 1496 1233 1504
rect 1247 1496 1313 1504
rect 1447 1496 1453 1504
rect 1467 1496 1593 1504
rect 2507 1496 3413 1504
rect 3427 1496 3453 1504
rect 3627 1496 4213 1504
rect 847 1476 1193 1484
rect 1207 1476 1413 1484
rect 1507 1476 1693 1484
rect 1707 1476 1793 1484
rect 207 1456 453 1464
rect 747 1456 853 1464
rect 887 1456 1553 1464
rect 3607 1456 3653 1464
rect 307 1436 373 1444
rect 387 1436 1033 1444
rect 1187 1436 1513 1444
rect 367 1416 413 1424
rect 827 1416 933 1424
rect 1447 1416 1533 1424
rect 4267 1416 4293 1424
rect 67 1396 73 1404
rect 87 1396 353 1404
rect 367 1396 433 1404
rect 1267 1396 1393 1404
rect 1407 1396 1413 1404
rect 1427 1396 1553 1404
rect 1747 1396 1833 1404
rect 1847 1396 1853 1404
rect 4187 1396 4293 1404
rect 107 1376 133 1384
rect 336 1376 393 1384
rect 236 1347 244 1373
rect 287 1356 324 1364
rect 67 1336 124 1344
rect 116 1327 124 1336
rect 187 1336 224 1344
rect 216 1324 224 1336
rect 256 1344 264 1353
rect 256 1336 284 1344
rect 216 1316 253 1324
rect 96 1304 104 1313
rect 96 1296 153 1304
rect 276 1304 284 1336
rect 316 1324 324 1356
rect 336 1347 344 1376
rect 407 1376 713 1384
rect 967 1376 1193 1384
rect 1487 1376 1524 1384
rect 776 1356 833 1364
rect 356 1327 364 1353
rect 376 1336 393 1344
rect 316 1316 344 1324
rect 336 1307 344 1316
rect 376 1307 384 1336
rect 427 1336 504 1344
rect 496 1327 504 1336
rect 696 1336 733 1344
rect 627 1316 644 1324
rect 187 1296 284 1304
rect 87 1276 133 1284
rect 147 1276 313 1284
rect 416 1284 424 1313
rect 496 1304 504 1313
rect 367 1276 424 1284
rect 476 1296 504 1304
rect 476 1264 484 1296
rect 516 1284 524 1313
rect 536 1304 544 1313
rect 636 1304 644 1316
rect 696 1324 704 1336
rect 667 1316 704 1324
rect 716 1304 724 1313
rect 536 1296 624 1304
rect 636 1296 724 1304
rect 616 1287 624 1296
rect 716 1287 724 1296
rect 776 1304 784 1356
rect 907 1356 973 1364
rect 1107 1356 1204 1364
rect 1027 1336 1033 1344
rect 1047 1336 1073 1344
rect 1127 1336 1173 1344
rect 1196 1344 1204 1356
rect 1227 1356 1373 1364
rect 1407 1356 1493 1364
rect 1516 1364 1524 1376
rect 1947 1376 2053 1384
rect 2067 1376 2093 1384
rect 3267 1376 3293 1384
rect 4187 1376 4393 1384
rect 1516 1356 1544 1364
rect 1196 1336 1224 1344
rect 796 1307 804 1333
rect 836 1307 844 1333
rect 916 1307 924 1333
rect 976 1324 984 1333
rect 947 1316 1093 1324
rect 1127 1316 1193 1324
rect 747 1296 784 1304
rect 1107 1296 1153 1304
rect 507 1276 524 1284
rect 567 1276 593 1284
rect 767 1276 813 1284
rect 867 1276 913 1284
rect 1216 1284 1224 1336
rect 1287 1336 1364 1344
rect 1276 1316 1333 1324
rect 1276 1304 1284 1316
rect 1356 1324 1364 1336
rect 1476 1336 1513 1344
rect 1356 1316 1433 1324
rect 1456 1307 1464 1333
rect 1267 1296 1284 1304
rect 1307 1296 1344 1304
rect 1007 1276 1224 1284
rect 1236 1276 1313 1284
rect 67 1256 484 1264
rect 607 1256 693 1264
rect 1007 1256 1053 1264
rect 1236 1264 1244 1276
rect 1336 1284 1344 1296
rect 1476 1284 1484 1336
rect 1536 1327 1544 1356
rect 1687 1356 1913 1364
rect 1927 1356 2184 1364
rect 1596 1336 1753 1344
rect 1596 1307 1604 1336
rect 1947 1336 1993 1344
rect 2007 1336 2024 1344
rect 1787 1316 1804 1324
rect 1616 1304 1624 1313
rect 1616 1296 1693 1304
rect 1796 1304 1804 1316
rect 1827 1316 1913 1324
rect 2016 1324 2024 1336
rect 2176 1327 2184 1356
rect 2456 1356 2653 1364
rect 2207 1336 2273 1344
rect 2367 1336 2433 1344
rect 2456 1344 2464 1356
rect 2987 1356 3173 1364
rect 3187 1356 3253 1364
rect 4147 1356 4213 1364
rect 4227 1356 4473 1364
rect 4647 1356 4673 1364
rect 4707 1356 4773 1364
rect 2447 1336 2464 1344
rect 2487 1336 2593 1344
rect 2727 1336 2813 1344
rect 3107 1336 3213 1344
rect 3747 1336 3853 1344
rect 3887 1336 3953 1344
rect 3967 1336 4733 1344
rect 2016 1316 2033 1324
rect 2047 1316 2153 1324
rect 1796 1296 1873 1304
rect 1996 1304 2004 1313
rect 1947 1296 2004 1304
rect 2196 1304 2204 1333
rect 2527 1316 2773 1324
rect 2827 1316 2993 1324
rect 3016 1316 3533 1324
rect 2167 1296 2204 1304
rect 2267 1296 2333 1304
rect 2607 1296 2633 1304
rect 2687 1296 2753 1304
rect 3016 1304 3024 1316
rect 3547 1316 3604 1324
rect 3596 1307 3604 1316
rect 3696 1316 3753 1324
rect 2847 1296 3024 1304
rect 3067 1296 3073 1304
rect 3087 1296 3113 1304
rect 1336 1276 1484 1284
rect 1507 1276 1653 1284
rect 1667 1276 1713 1284
rect 1807 1276 1893 1284
rect 1987 1276 2073 1284
rect 2087 1276 2133 1284
rect 2467 1276 2493 1284
rect 2987 1276 3393 1284
rect 3476 1284 3484 1293
rect 3616 1287 3624 1313
rect 3696 1304 3704 1316
rect 3767 1316 4053 1324
rect 4107 1316 4153 1324
rect 4347 1316 4393 1324
rect 4496 1316 4533 1324
rect 3647 1296 3704 1304
rect 3727 1296 3813 1304
rect 3947 1296 4073 1304
rect 4387 1296 4413 1304
rect 3476 1276 3553 1284
rect 3567 1276 3593 1284
rect 3647 1276 3673 1284
rect 3707 1276 3793 1284
rect 4436 1284 4444 1313
rect 4496 1307 4504 1316
rect 4727 1316 4753 1324
rect 4787 1316 4824 1324
rect 4676 1304 4684 1313
rect 4567 1296 4684 1304
rect 4436 1276 4513 1284
rect 4587 1276 4653 1284
rect 1067 1256 1244 1264
rect 1267 1256 1333 1264
rect 1387 1256 1533 1264
rect 1567 1256 1693 1264
rect 1847 1256 1933 1264
rect 1967 1256 2093 1264
rect 2947 1256 3193 1264
rect 3247 1256 3873 1264
rect 4467 1256 4593 1264
rect 447 1236 573 1244
rect 647 1236 853 1244
rect 887 1236 1193 1244
rect 1587 1236 2013 1244
rect 2147 1236 2213 1244
rect 2807 1236 3353 1244
rect 3407 1236 3613 1244
rect 3956 1236 4033 1244
rect 287 1216 453 1224
rect 467 1216 513 1224
rect 587 1216 713 1224
rect 807 1216 853 1224
rect 907 1216 1024 1224
rect 307 1196 553 1204
rect 627 1196 713 1204
rect 807 1196 993 1204
rect 1016 1204 1024 1216
rect 1207 1216 1393 1224
rect 1867 1216 2013 1224
rect 3956 1224 3964 1236
rect 3467 1216 3964 1224
rect 1016 1196 1053 1204
rect 1147 1196 1353 1204
rect 1627 1196 1773 1204
rect 2707 1196 3273 1204
rect 3287 1196 3373 1204
rect 3947 1196 4013 1204
rect -4 1176 213 1184
rect -4 1124 4 1176
rect 307 1176 333 1184
rect 387 1176 593 1184
rect 627 1176 653 1184
rect 747 1176 1033 1184
rect 1187 1176 1213 1184
rect 1587 1176 1633 1184
rect 2647 1176 2853 1184
rect 3387 1176 4273 1184
rect 167 1156 373 1164
rect 407 1156 413 1164
rect 427 1156 653 1164
rect 847 1156 893 1164
rect 987 1156 1093 1164
rect 1147 1156 1193 1164
rect 1527 1156 1693 1164
rect 2687 1156 2873 1164
rect 2907 1156 2973 1164
rect 3147 1156 3473 1164
rect 4447 1156 4573 1164
rect 27 1136 93 1144
rect 107 1136 113 1144
rect 156 1136 204 1144
rect -4 1116 13 1124
rect 47 1116 84 1124
rect 76 1107 84 1116
rect 87 1096 133 1104
rect 36 1084 44 1093
rect 36 1076 93 1084
rect 156 1084 164 1136
rect 107 1076 164 1084
rect 176 1067 184 1113
rect 196 1104 204 1136
rect 247 1136 333 1144
rect 447 1136 533 1144
rect 567 1136 584 1144
rect 227 1116 253 1124
rect 267 1116 293 1124
rect 356 1124 364 1133
rect 356 1116 373 1124
rect 427 1116 564 1124
rect 556 1107 564 1116
rect 196 1096 253 1104
rect 376 1096 433 1104
rect 376 1084 384 1096
rect 467 1096 513 1104
rect 287 1076 384 1084
rect 456 1084 464 1093
rect 576 1087 584 1136
rect 847 1136 1033 1144
rect 1056 1136 1113 1144
rect 856 1116 933 1124
rect 736 1087 744 1113
rect 776 1087 784 1113
rect 407 1076 464 1084
rect 487 1076 533 1084
rect 687 1076 733 1084
rect 207 1056 253 1064
rect 267 1056 353 1064
rect 507 1056 533 1064
rect 816 1064 824 1113
rect 856 1107 864 1116
rect 1056 1107 1064 1136
rect 1127 1136 1233 1144
rect 1307 1136 1353 1144
rect 1367 1136 1613 1144
rect 1647 1136 1673 1144
rect 1707 1136 1793 1144
rect 1867 1136 2053 1144
rect 2227 1136 2353 1144
rect 2627 1136 2693 1144
rect 3007 1136 3173 1144
rect 3187 1136 3213 1144
rect 3227 1136 3333 1144
rect 3827 1136 3853 1144
rect 3907 1136 4133 1144
rect 4187 1136 4393 1144
rect 4567 1136 4753 1144
rect 1127 1116 1293 1124
rect 1216 1087 1224 1116
rect 1447 1116 1473 1124
rect 1487 1116 1553 1124
rect 1687 1116 1753 1124
rect 1767 1116 1873 1124
rect 1936 1116 2133 1124
rect 1247 1096 1364 1104
rect 1356 1087 1364 1096
rect 1376 1087 1384 1113
rect 1416 1104 1424 1113
rect 1416 1096 1493 1104
rect 1567 1096 1624 1104
rect 1616 1087 1624 1096
rect 1827 1096 1893 1104
rect 1936 1104 1944 1116
rect 2407 1116 2593 1124
rect 2656 1116 2733 1124
rect 2656 1107 2664 1116
rect 2747 1116 2793 1124
rect 2987 1116 3013 1124
rect 3267 1116 3573 1124
rect 3587 1116 3593 1124
rect 3607 1116 3873 1124
rect 3927 1116 4013 1124
rect 4027 1116 4293 1124
rect 4307 1116 4333 1124
rect 4347 1116 4353 1124
rect 4376 1116 4444 1124
rect 4376 1107 4384 1116
rect 1916 1096 1944 1104
rect 967 1076 1153 1084
rect 1427 1076 1453 1084
rect 1467 1076 1473 1084
rect 1716 1084 1724 1093
rect 1916 1087 1924 1096
rect 2127 1096 2153 1104
rect 2207 1096 2373 1104
rect 2387 1096 2453 1104
rect 2547 1096 2613 1104
rect 3047 1096 3113 1104
rect 3427 1096 3493 1104
rect 3507 1096 3693 1104
rect 3847 1096 3853 1104
rect 3867 1096 3893 1104
rect 3987 1096 4033 1104
rect 4307 1096 4364 1104
rect 1667 1076 1724 1084
rect 1747 1076 1873 1084
rect 2087 1076 2173 1084
rect 2187 1076 2273 1084
rect 2287 1076 2513 1084
rect 2567 1076 2653 1084
rect 4067 1076 4193 1084
rect 4207 1076 4273 1084
rect 4356 1084 4364 1096
rect 4436 1104 4444 1116
rect 4507 1116 4564 1124
rect 4556 1107 4564 1116
rect 4647 1116 4673 1124
rect 4707 1116 4733 1124
rect 4436 1096 4493 1104
rect 4576 1096 4593 1104
rect 4416 1084 4424 1093
rect 4356 1076 4424 1084
rect 4447 1076 4473 1084
rect 4576 1084 4584 1096
rect 4567 1076 4584 1084
rect 4667 1076 4684 1084
rect 4676 1067 4684 1076
rect 816 1056 873 1064
rect 907 1056 1313 1064
rect 1327 1056 1393 1064
rect 1627 1056 1793 1064
rect 1847 1056 1933 1064
rect 2047 1056 2253 1064
rect 2267 1056 2313 1064
rect 2927 1056 2993 1064
rect 567 1036 1573 1044
rect 1587 1036 1753 1044
rect 1827 1036 1953 1044
rect 4527 1036 4693 1044
rect 647 1016 773 1024
rect 787 1016 813 1024
rect 1307 1016 1624 1024
rect 787 996 1533 1004
rect 1616 1004 1624 1016
rect 1647 1016 1893 1024
rect 1907 1016 2013 1024
rect 1616 996 1653 1004
rect 847 976 893 984
rect 1167 976 1433 984
rect 1507 976 1753 984
rect 1807 976 2513 984
rect 3667 976 3913 984
rect 3927 976 3953 984
rect 1007 956 1073 964
rect 1187 956 1253 964
rect 1267 956 1813 964
rect 2507 956 2553 964
rect 27 936 893 944
rect 1087 936 1193 944
rect 1547 936 1653 944
rect 1787 936 2153 944
rect 527 916 753 924
rect 767 916 813 924
rect 1027 916 1113 924
rect 1207 916 1313 924
rect 1367 916 1433 924
rect 1496 916 1604 924
rect 507 896 573 904
rect 867 896 913 904
rect 927 896 1213 904
rect 1407 896 1453 904
rect 1496 904 1504 916
rect 1467 896 1504 904
rect 1596 904 1604 916
rect 1627 916 1833 924
rect 4507 916 4613 924
rect 4667 916 4753 924
rect 1596 896 1633 904
rect 1667 896 1933 904
rect 4567 896 4753 904
rect 87 876 293 884
rect 427 876 693 884
rect 1056 876 1073 884
rect 1056 867 1064 876
rect 1227 876 1273 884
rect 1387 876 1553 884
rect 1536 867 1544 876
rect 1607 876 1733 884
rect 1747 876 1833 884
rect 1947 876 1993 884
rect 2007 876 2413 884
rect 4627 876 4733 884
rect 236 856 253 864
rect 236 827 244 856
rect 276 856 364 864
rect 276 844 284 856
rect 267 836 284 844
rect 127 816 133 824
rect 147 816 193 824
rect 27 796 153 804
rect 336 804 344 833
rect 356 827 364 856
rect 387 856 453 864
rect 587 856 653 864
rect 707 856 733 864
rect 847 856 864 864
rect 396 836 493 844
rect 396 827 404 836
rect 607 836 644 844
rect 636 807 644 836
rect 707 836 844 844
rect 836 827 844 836
rect 856 827 864 856
rect 907 856 944 864
rect 936 844 944 856
rect 967 856 973 864
rect 987 856 1013 864
rect 1127 856 1333 864
rect 1347 856 1373 864
rect 1396 856 1473 864
rect 936 836 1053 844
rect 1096 827 1104 853
rect 1207 836 1253 844
rect 1396 844 1404 856
rect 1587 856 1753 864
rect 1767 856 1873 864
rect 1987 856 2353 864
rect 2367 856 2444 864
rect 2436 847 2444 856
rect 2507 856 2544 864
rect 1347 836 1404 844
rect 1427 836 1553 844
rect 1567 836 1673 844
rect 1756 836 2053 844
rect 696 816 753 824
rect 167 796 433 804
rect 447 796 493 804
rect 696 804 704 816
rect 907 816 973 824
rect 1296 824 1304 833
rect 1756 827 1764 836
rect 2147 836 2193 844
rect 2327 836 2393 844
rect 2536 844 2544 856
rect 2567 856 2753 864
rect 2807 856 2893 864
rect 2907 856 2933 864
rect 3367 856 3393 864
rect 3647 856 3713 864
rect 3947 856 4013 864
rect 2536 836 2573 844
rect 2607 836 2633 844
rect 2787 836 2853 844
rect 3087 836 3233 844
rect 1296 816 1553 824
rect 1607 816 1713 824
rect 1787 816 1813 824
rect 1896 816 2173 824
rect 687 796 704 804
rect 727 796 933 804
rect 1107 796 1353 804
rect 1727 796 1793 804
rect 1896 804 1904 816
rect 2227 816 2273 824
rect 2676 824 2684 833
rect 2627 816 2684 824
rect 2707 816 2833 824
rect 2956 824 2964 833
rect 2927 816 3044 824
rect 1836 796 1904 804
rect 187 776 293 784
rect 707 776 873 784
rect 1087 776 1293 784
rect 1307 776 1493 784
rect 1836 784 1844 796
rect 1927 796 1953 804
rect 2027 796 2173 804
rect 2247 796 2293 804
rect 2587 796 2653 804
rect 2987 796 3013 804
rect 3036 804 3044 816
rect 3067 816 3164 824
rect 3156 807 3164 816
rect 3316 824 3324 853
rect 3347 836 3373 844
rect 4036 844 4044 853
rect 3987 836 4044 844
rect 3267 816 3324 824
rect 3487 816 3533 824
rect 3607 816 3633 824
rect 3807 816 3993 824
rect 4087 816 4253 824
rect 4267 816 4313 824
rect 4467 816 4633 824
rect 3036 796 3093 804
rect 3416 804 3424 813
rect 4676 807 4684 853
rect 3167 796 3424 804
rect 3507 796 3713 804
rect 3867 796 4113 804
rect 4127 796 4153 804
rect 4167 796 4173 804
rect 4187 796 4413 804
rect 4427 796 4633 804
rect 1727 776 1844 784
rect 1867 776 1933 784
rect 1947 776 1993 784
rect 2067 776 2253 784
rect 3087 776 3113 784
rect 3147 776 3193 784
rect 3947 776 4073 784
rect 4387 776 4693 784
rect 607 756 653 764
rect 667 756 733 764
rect 1047 756 1133 764
rect 1287 756 1393 764
rect 1427 756 1613 764
rect 1747 756 1833 764
rect 2007 756 2193 764
rect 2207 756 2433 764
rect 3007 756 3073 764
rect 3347 756 3393 764
rect 4207 756 4453 764
rect 487 736 533 744
rect 547 736 553 744
rect 567 736 773 744
rect 1247 736 1433 744
rect 1487 736 1753 744
rect 1987 736 2133 744
rect 2287 736 2573 744
rect 547 716 993 724
rect 1247 716 1684 724
rect 227 696 253 704
rect 267 696 393 704
rect 427 696 613 704
rect 827 696 893 704
rect 967 696 1193 704
rect 1327 696 1333 704
rect 1347 696 1493 704
rect 1507 696 1653 704
rect 1676 704 1684 716
rect 1707 716 1953 724
rect 1967 716 2033 724
rect 2047 716 2533 724
rect 2927 716 2953 724
rect 2967 716 3493 724
rect 3787 716 4213 724
rect 1676 696 2053 704
rect 2107 696 2373 704
rect 2387 696 2453 704
rect 167 676 313 684
rect 327 676 353 684
rect 447 676 673 684
rect 807 676 913 684
rect 1027 676 1113 684
rect 1287 676 1353 684
rect 1447 676 1533 684
rect 1607 676 1733 684
rect 1887 676 2233 684
rect 2347 676 2373 684
rect 2387 676 2473 684
rect 3367 676 3513 684
rect 3687 676 3833 684
rect 3847 676 3933 684
rect 3947 676 4033 684
rect 4047 676 4393 684
rect 4407 676 4493 684
rect 67 656 104 664
rect 96 624 104 656
rect 147 656 164 664
rect 156 627 164 656
rect 207 656 273 664
rect 316 656 373 664
rect 196 627 204 653
rect 247 636 273 644
rect 316 627 324 656
rect 467 656 524 664
rect 367 636 493 644
rect 516 644 524 656
rect 627 656 833 664
rect 887 656 993 664
rect 1007 656 1033 664
rect 1067 656 1084 664
rect 516 636 573 644
rect 596 636 633 644
rect 96 616 133 624
rect 347 616 393 624
rect 596 624 604 636
rect 656 636 713 644
rect 487 616 504 624
rect 496 607 504 616
rect 516 616 604 624
rect 187 596 213 604
rect 227 596 293 604
rect 307 596 373 604
rect 516 587 524 616
rect 656 624 664 636
rect 827 636 853 644
rect 867 636 884 644
rect 647 616 664 624
rect 876 607 884 636
rect 1027 636 1053 644
rect 1076 627 1084 656
rect 1467 656 1513 664
rect 1576 656 1593 664
rect 1107 636 1133 644
rect 1387 636 1413 644
rect 1576 644 1584 656
rect 1667 656 1713 664
rect 1787 656 1813 664
rect 2096 656 2113 664
rect 2016 644 2024 653
rect 2096 644 2104 656
rect 2327 656 2333 664
rect 2347 656 2413 664
rect 2467 656 2513 664
rect 3047 656 3193 664
rect 3207 656 3213 664
rect 3247 656 3273 664
rect 3287 656 3393 664
rect 3467 656 3493 664
rect 3507 656 3573 664
rect 3827 656 4013 664
rect 1476 636 1584 644
rect 1736 636 2024 644
rect 2076 636 2104 644
rect 907 616 933 624
rect 987 616 1013 624
rect 1127 616 1173 624
rect 1227 616 1253 624
rect 1476 624 1484 636
rect 1307 616 1484 624
rect 1736 624 1744 636
rect 1607 616 1744 624
rect 1767 616 1844 624
rect 1836 607 1844 616
rect 2076 624 2084 636
rect 2127 636 2213 644
rect 2267 636 2304 644
rect 2296 627 2304 636
rect 2407 636 2473 644
rect 2676 627 2684 653
rect 2707 636 2773 644
rect 2787 636 2933 644
rect 3187 636 3253 644
rect 3307 636 3413 644
rect 3547 636 3673 644
rect 3887 636 3913 644
rect 3967 636 4033 644
rect 4107 636 4153 644
rect 4667 636 4673 644
rect 4687 636 4713 644
rect 2007 616 2084 624
rect 2107 616 2144 624
rect 787 596 853 604
rect 1087 596 1373 604
rect 1467 596 1573 604
rect 1727 596 1753 604
rect 1987 596 2113 604
rect 2136 604 2144 616
rect 2307 616 2353 624
rect 2376 616 2453 624
rect 2136 596 2153 604
rect 287 576 513 584
rect 547 576 893 584
rect 1427 576 1673 584
rect 1756 584 1764 593
rect 2176 587 2184 613
rect 2207 596 2273 604
rect 2376 604 2384 616
rect 2487 616 2513 624
rect 2696 616 2733 624
rect 2307 596 2384 604
rect 2507 596 2553 604
rect 2696 604 2704 616
rect 3107 616 3153 624
rect 3167 616 3273 624
rect 3307 616 3373 624
rect 3467 616 3513 624
rect 3567 616 3813 624
rect 3907 616 3973 624
rect 4247 616 4273 624
rect 4367 616 4433 624
rect 2667 596 2704 604
rect 3067 596 3233 604
rect 4007 596 4033 604
rect 4227 596 4253 604
rect 1687 576 1764 584
rect 1787 576 1853 584
rect 1907 576 2164 584
rect 567 556 2093 564
rect 2156 564 2164 576
rect 2456 584 2464 593
rect 2187 576 2464 584
rect 2716 564 2724 593
rect 3187 576 3213 584
rect 3927 576 4093 584
rect 2156 556 2724 564
rect 707 536 773 544
rect 1127 536 1153 544
rect 1167 536 1493 544
rect 1527 536 1653 544
rect 1676 536 1813 544
rect 327 516 473 524
rect 1367 516 1533 524
rect 1567 516 1593 524
rect 1676 524 1684 536
rect 1827 536 2013 544
rect 2047 536 2173 544
rect 2687 536 2733 544
rect 3807 536 3993 544
rect 1647 516 1684 524
rect 1707 516 1833 524
rect 2067 516 2133 524
rect 4487 516 4693 524
rect 367 496 433 504
rect 527 496 613 504
rect 627 496 1073 504
rect 1227 496 1733 504
rect 1847 496 2413 504
rect 447 476 493 484
rect 1727 476 1773 484
rect 1807 476 1993 484
rect 2147 476 2173 484
rect 2187 476 2293 484
rect 327 456 513 464
rect 527 456 873 464
rect 1407 456 1873 464
rect 1927 456 2193 464
rect 407 436 633 444
rect 987 436 1273 444
rect 1367 436 1593 444
rect 1607 436 1853 444
rect 1927 436 2273 444
rect 247 416 333 424
rect 547 416 593 424
rect 887 416 993 424
rect 1147 416 1353 424
rect 1387 416 1693 424
rect 1727 416 1893 424
rect 2047 416 2113 424
rect 2127 416 2413 424
rect 2567 416 2633 424
rect 2647 416 2873 424
rect 3487 416 3893 424
rect 3907 416 4293 424
rect 4307 416 4473 424
rect 4487 416 4533 424
rect 107 396 433 404
rect 467 396 653 404
rect 707 396 853 404
rect 867 396 933 404
rect 947 396 1173 404
rect 1467 396 1633 404
rect 1667 396 1804 404
rect 167 376 193 384
rect 316 376 353 384
rect 227 356 253 364
rect 316 347 324 376
rect 387 376 453 384
rect 507 376 724 384
rect 407 356 593 364
rect 716 347 724 376
rect 907 376 1004 384
rect 836 364 844 373
rect 836 356 953 364
rect 107 336 173 344
rect 187 336 293 344
rect 427 336 713 344
rect 87 316 253 324
rect 267 316 353 324
rect 447 316 473 324
rect 527 316 633 324
rect 776 324 784 353
rect 996 344 1004 376
rect 1127 376 1244 384
rect 1027 356 1133 364
rect 1236 347 1244 376
rect 1287 376 1333 384
rect 1587 376 1664 384
rect 1256 347 1264 373
rect 1327 356 1353 364
rect 1407 356 1424 364
rect 1416 347 1424 356
rect 1456 356 1533 364
rect 827 336 964 344
rect 996 336 1153 344
rect 707 316 784 324
rect 807 316 913 324
rect 956 324 964 336
rect 1456 327 1464 356
rect 1556 344 1564 373
rect 1487 336 1564 344
rect 956 316 993 324
rect 1067 316 1113 324
rect 1187 316 1413 324
rect 1636 324 1644 353
rect 1487 316 1644 324
rect 1656 324 1664 376
rect 1796 384 1804 396
rect 1827 396 1913 404
rect 1967 396 2333 404
rect 2587 396 2693 404
rect 2767 396 3613 404
rect 3647 396 3793 404
rect 4287 396 4353 404
rect 1687 376 1784 384
rect 1796 376 1824 384
rect 1687 356 1713 364
rect 1727 356 1753 364
rect 1776 344 1784 376
rect 1816 347 1824 376
rect 1947 376 1993 384
rect 2107 376 2213 384
rect 2347 376 2444 384
rect 1887 356 2013 364
rect 2027 356 2053 364
rect 1747 336 1784 344
rect 1847 336 1913 344
rect 2076 344 2084 373
rect 2436 367 2444 376
rect 2507 376 2533 384
rect 2556 376 2733 384
rect 2147 356 2193 364
rect 2247 356 2384 364
rect 2067 336 2273 344
rect 2327 336 2353 344
rect 2376 344 2384 356
rect 2556 364 2564 376
rect 2676 367 2684 376
rect 2867 376 2893 384
rect 2947 376 3013 384
rect 3027 376 3113 384
rect 3316 376 3353 384
rect 3316 367 3324 376
rect 3407 376 3473 384
rect 4327 376 4373 384
rect 2456 356 2564 364
rect 2376 336 2433 344
rect 1656 316 1673 324
rect 1707 316 1853 324
rect 2027 316 2213 324
rect 2456 324 2464 356
rect 2587 356 2633 364
rect 2696 356 2773 364
rect 2696 344 2704 356
rect 2927 356 3073 364
rect 3756 364 3764 373
rect 3707 356 3764 364
rect 3787 356 3833 364
rect 4087 356 4333 364
rect 4447 356 4493 364
rect 2487 336 2704 344
rect 2767 336 2793 344
rect 2847 336 2873 344
rect 3147 336 3173 344
rect 3356 344 3364 353
rect 3247 336 3364 344
rect 3436 344 3444 353
rect 3436 336 3513 344
rect 3627 336 3853 344
rect 4087 336 4113 344
rect 4267 336 4393 344
rect 2387 316 2464 324
rect 2667 316 2713 324
rect 2827 316 2853 324
rect 3067 316 3413 324
rect 3467 316 3533 324
rect 3547 316 3593 324
rect 3607 316 3653 324
rect 4047 316 4133 324
rect 4496 324 4504 353
rect 4487 316 4504 324
rect 487 296 753 304
rect 827 296 1033 304
rect 1047 296 1133 304
rect 1267 296 1493 304
rect 1507 296 1693 304
rect 1767 296 1953 304
rect 2007 296 2033 304
rect 2147 296 2253 304
rect 2267 296 2393 304
rect 2547 296 2973 304
rect 3107 296 3353 304
rect 3507 296 3573 304
rect 3587 296 3733 304
rect 3747 296 3933 304
rect 3987 296 4113 304
rect 4427 296 4673 304
rect 367 276 953 284
rect 1207 276 1333 284
rect 1347 276 1433 284
rect 1447 276 1533 284
rect 1607 276 1793 284
rect 2207 276 2253 284
rect 3207 276 3513 284
rect 3887 276 4193 284
rect 367 256 553 264
rect 927 256 1373 264
rect 1407 256 1473 264
rect 1587 256 1653 264
rect 1667 256 1773 264
rect 1787 256 1873 264
rect 1987 256 2393 264
rect 2407 256 2653 264
rect 2667 256 2693 264
rect 3287 256 3573 264
rect 3927 256 3973 264
rect 3987 256 4033 264
rect 427 236 733 244
rect 907 236 1273 244
rect 1287 236 1373 244
rect 1427 236 1633 244
rect 1707 236 2073 244
rect 2967 236 3013 244
rect 3347 236 3733 244
rect 687 216 813 224
rect 867 216 893 224
rect 1027 216 1093 224
rect 1127 216 2013 224
rect 2147 216 2173 224
rect 2187 216 2193 224
rect 2207 216 2453 224
rect 3087 216 3153 224
rect 3967 216 4373 224
rect 47 196 133 204
rect 247 196 553 204
rect 627 196 853 204
rect 967 196 1033 204
rect 1087 196 1213 204
rect 1307 196 1533 204
rect 1627 196 1773 204
rect 2107 196 2153 204
rect 2187 196 2253 204
rect 2367 196 2413 204
rect 2567 196 2773 204
rect 3047 196 3193 204
rect 3207 196 4513 204
rect 87 176 113 184
rect 267 176 313 184
rect 447 176 473 184
rect 487 176 533 184
rect 547 176 633 184
rect 807 176 973 184
rect 1007 176 1313 184
rect 1447 176 1493 184
rect 1527 176 1673 184
rect 1707 176 1733 184
rect 1967 176 2053 184
rect 2087 176 2353 184
rect 2607 176 2853 184
rect 3047 176 3393 184
rect 3407 176 3693 184
rect 3807 176 3833 184
rect 3847 176 3993 184
rect 4027 176 4173 184
rect 4207 176 4333 184
rect 4427 176 4453 184
rect 4467 176 4493 184
rect 4527 176 4613 184
rect 107 156 164 164
rect 156 147 164 156
rect 187 156 293 164
rect 307 156 313 164
rect 336 147 344 173
rect 387 156 493 164
rect 507 156 593 164
rect 616 156 733 164
rect 87 136 113 144
rect 287 136 333 144
rect 467 136 513 144
rect 616 144 624 156
rect 756 147 764 173
rect 776 164 784 173
rect 776 156 864 164
rect 567 136 624 144
rect 807 136 833 144
rect 856 144 864 156
rect 887 156 913 164
rect 936 156 1093 164
rect 936 147 944 156
rect 1107 156 1333 164
rect 1447 156 1553 164
rect 1596 156 1753 164
rect 856 136 904 144
rect 516 124 524 133
rect 47 116 524 124
rect 516 104 524 116
rect 607 116 653 124
rect 667 116 873 124
rect 896 124 904 136
rect 987 136 1053 144
rect 1067 136 1113 144
rect 1156 136 1193 144
rect 896 116 993 124
rect 1156 124 1164 136
rect 1207 136 1233 144
rect 1336 136 1433 144
rect 1007 116 1164 124
rect 1236 116 1253 124
rect 516 96 613 104
rect 1236 104 1244 116
rect 1336 124 1344 136
rect 1487 136 1533 144
rect 1307 116 1344 124
rect 1576 124 1584 133
rect 1596 127 1604 156
rect 1927 156 1973 164
rect 2027 156 2213 164
rect 2327 156 2593 164
rect 2416 147 2424 156
rect 2787 156 2824 164
rect 1627 136 1673 144
rect 1707 136 1733 144
rect 1936 136 2173 144
rect 1527 116 1584 124
rect 1647 116 1713 124
rect 1727 116 1753 124
rect 1827 116 1893 124
rect 1936 124 1944 136
rect 2207 136 2333 144
rect 2587 136 2713 144
rect 2727 136 2753 144
rect 2816 144 2824 156
rect 3087 156 3113 164
rect 3287 156 3473 164
rect 3487 156 3533 164
rect 3587 156 3613 164
rect 3827 156 3873 164
rect 3887 156 3893 164
rect 3907 156 3993 164
rect 4016 156 4073 164
rect 2816 136 2873 144
rect 3147 136 3233 144
rect 4016 144 4024 156
rect 4487 156 4533 164
rect 3807 136 4024 144
rect 4216 144 4224 153
rect 4067 136 4253 144
rect 4307 136 4433 144
rect 4587 136 4644 144
rect 1927 116 1944 124
rect 2267 116 2533 124
rect 2547 116 2613 124
rect 1356 104 1364 113
rect 847 96 1364 104
rect 1407 96 1693 104
rect 1807 96 1993 104
rect 2247 96 2473 104
rect 2796 104 2804 133
rect 3927 116 3973 124
rect 4636 124 4644 136
rect 4667 136 4753 144
rect 4636 116 4693 124
rect 2487 96 2804 104
rect 4447 96 4733 104
rect 987 76 1473 84
rect 1847 76 1913 84
rect 2067 76 2293 84
rect 2747 76 2813 84
rect 1227 56 1513 64
rect 1767 56 2113 64
rect 867 36 1873 44
rect 1887 36 1933 44
rect 1327 16 1973 24
rect 2127 16 2153 24
<< m1p >>
rect 4 4562 4776 4578
rect 4 4322 4776 4338
rect 4 4082 4736 4098
rect 4 3842 4776 3858
rect 4 3602 4736 3618
rect 4 3362 4776 3378
rect 4 3122 4776 3138
rect 4 2882 4776 2898
rect 4 2642 4736 2658
rect 4 2402 4776 2418
rect 4 2162 4776 2178
rect 4 1922 4776 1938
rect 4 1682 4776 1698
rect 4 1442 4776 1458
rect 4 1202 4776 1218
rect 4 962 4776 978
rect 4 722 4756 738
rect 4 482 4776 498
rect 4 242 4776 258
rect 4 2 4776 18
<< m2p >>
rect 73 4493 87 4507
rect 433 4493 447 4507
rect 1113 4493 1127 4507
rect 1313 4493 1327 4507
rect 1553 4493 1567 4507
rect 1773 4493 1787 4507
rect 1813 4493 1827 4507
rect 1913 4493 1927 4507
rect 1953 4493 1967 4507
rect 2053 4493 2067 4507
rect 2113 4493 2127 4507
rect 2393 4493 2407 4507
rect 2513 4493 2527 4507
rect 2993 4493 3007 4507
rect 3153 4493 3167 4507
rect 3333 4493 3347 4507
rect 3413 4493 3427 4507
rect 4213 4493 4227 4507
rect 33 4473 47 4487
rect 473 4473 487 4487
rect 513 4473 527 4487
rect 553 4473 567 4487
rect 613 4473 627 4487
rect 653 4473 667 4487
rect 1153 4473 1167 4487
rect 1293 4473 1307 4487
rect 1333 4473 1347 4487
rect 1393 4473 1407 4487
rect 1433 4473 1447 4487
rect 1533 4473 1547 4487
rect 1573 4473 1587 4487
rect 1733 4473 1747 4487
rect 1993 4473 2007 4487
rect 2033 4473 2047 4487
rect 2073 4473 2087 4487
rect 2173 4473 2187 4487
rect 2213 4473 2227 4487
rect 2293 4473 2307 4487
rect 2333 4473 2347 4487
rect 2373 4473 2387 4487
rect 2413 4473 2427 4487
rect 2553 4473 2567 4487
rect 2613 4473 2627 4487
rect 2653 4473 2667 4487
rect 2693 4473 2707 4487
rect 2793 4473 2807 4487
rect 2833 4473 2847 4487
rect 2913 4473 2927 4487
rect 3053 4473 3067 4487
rect 3093 4473 3107 4487
rect 3133 4473 3147 4487
rect 3173 4473 3187 4487
rect 3233 4473 3247 4487
rect 3273 4473 3287 4487
rect 3313 4473 3327 4487
rect 3353 4473 3367 4487
rect 3453 4473 3467 4487
rect 3533 4473 3547 4487
rect 3573 4473 3587 4487
rect 3673 4473 3687 4487
rect 3713 4473 3727 4487
rect 4073 4473 4087 4487
rect 4113 4473 4127 4487
rect 4273 4473 4287 4487
rect 4313 4473 4327 4487
rect 4393 4473 4407 4487
rect 4473 4473 4487 4487
rect 4513 4473 4527 4487
rect 4613 4473 4627 4487
rect 4653 4473 4667 4487
rect 53 4453 67 4467
rect 93 4453 107 4467
rect 153 4453 167 4467
rect 193 4453 207 4467
rect 213 4453 227 4467
rect 253 4453 267 4467
rect 353 4453 367 4467
rect 393 4453 407 4467
rect 413 4453 427 4467
rect 453 4453 467 4467
rect 533 4453 547 4467
rect 573 4453 587 4467
rect 633 4453 647 4467
rect 673 4453 687 4467
rect 753 4453 767 4467
rect 793 4453 807 4467
rect 813 4453 827 4467
rect 853 4453 867 4467
rect 933 4453 947 4467
rect 993 4453 1007 4467
rect 1033 4453 1047 4467
rect 1093 4453 1107 4467
rect 1133 4453 1147 4467
rect 1233 4453 1247 4467
rect 1373 4453 1387 4467
rect 1413 4453 1427 4467
rect 1493 4453 1507 4467
rect 1613 4453 1627 4467
rect 1653 4453 1667 4467
rect 1753 4453 1767 4467
rect 1793 4453 1807 4467
rect 1833 4453 1847 4467
rect 1893 4453 1907 4467
rect 1933 4453 1947 4467
rect 1973 4453 1987 4467
rect 2133 4453 2147 4467
rect 2193 4453 2207 4467
rect 2233 4453 2247 4467
rect 2313 4453 2327 4467
rect 2353 4453 2367 4467
rect 2453 4453 2467 4467
rect 2493 4453 2507 4467
rect 2533 4453 2547 4467
rect 2633 4453 2647 4467
rect 2673 4453 2687 4467
rect 2973 4453 2987 4467
rect 3033 4453 3047 4467
rect 3073 4453 3087 4467
rect 3213 4453 3227 4467
rect 3253 4453 3267 4467
rect 3393 4453 3407 4467
rect 3693 4453 3707 4467
rect 3733 4453 3747 4467
rect 3793 4453 3807 4467
rect 3873 4453 3887 4467
rect 4013 4453 4027 4467
rect 4153 4453 4167 4467
rect 4233 4453 4247 4467
rect 4293 4453 4307 4467
rect 4333 4453 4347 4467
rect 4713 4453 4727 4467
rect 133 4433 147 4447
rect 173 4433 187 4447
rect 233 4433 247 4447
rect 273 4433 287 4447
rect 333 4433 347 4447
rect 373 4433 387 4447
rect 733 4433 747 4447
rect 773 4433 787 4447
rect 833 4433 847 4447
rect 873 4433 887 4447
rect 913 4433 927 4447
rect 953 4433 967 4447
rect 1013 4433 1027 4447
rect 1053 4433 1067 4447
rect 1213 4433 1227 4447
rect 1253 4433 1267 4447
rect 1473 4433 1487 4447
rect 1513 4433 1527 4447
rect 1633 4433 1647 4447
rect 1673 4433 1687 4447
rect 3773 4433 3787 4447
rect 3813 4433 3827 4447
rect 4133 4433 4147 4447
rect 4173 4433 4187 4447
rect 4693 4433 4707 4447
rect 4733 4433 4747 4447
rect 33 4213 47 4227
rect 73 4213 87 4227
rect 213 4213 227 4227
rect 253 4213 267 4227
rect 793 4213 807 4227
rect 833 4213 847 4227
rect 1013 4213 1027 4227
rect 1053 4213 1067 4227
rect 1113 4213 1127 4227
rect 1153 4213 1167 4227
rect 1213 4213 1227 4227
rect 1253 4213 1267 4227
rect 1293 4213 1307 4227
rect 1333 4213 1347 4227
rect 1393 4213 1407 4227
rect 1433 4213 1447 4227
rect 1473 4213 1487 4227
rect 1513 4213 1527 4227
rect 1833 4213 1847 4227
rect 1873 4213 1887 4227
rect 1973 4213 1987 4227
rect 2013 4213 2027 4227
rect 2073 4213 2087 4227
rect 2113 4213 2127 4227
rect 3093 4213 3107 4227
rect 3133 4213 3147 4227
rect 3193 4213 3207 4227
rect 3233 4213 3247 4227
rect 3273 4213 3287 4227
rect 3313 4213 3327 4227
rect 3673 4213 3687 4227
rect 3713 4213 3727 4227
rect 53 4193 67 4207
rect 93 4193 107 4207
rect 133 4193 147 4207
rect 233 4193 247 4207
rect 373 4193 387 4207
rect 413 4193 427 4207
rect 473 4193 487 4207
rect 513 4193 527 4207
rect 573 4193 587 4207
rect 653 4193 667 4207
rect 693 4193 707 4207
rect 733 4193 747 4207
rect 773 4193 787 4207
rect 813 4193 827 4207
rect 913 4193 927 4207
rect 953 4193 967 4207
rect 1033 4193 1047 4207
rect 1073 4193 1087 4207
rect 1093 4193 1107 4207
rect 1133 4193 1147 4207
rect 1233 4193 1247 4207
rect 1313 4193 1327 4207
rect 1353 4193 1367 4207
rect 1413 4193 1427 4207
rect 1453 4193 1467 4207
rect 1493 4193 1507 4207
rect 1733 4193 1747 4207
rect 1773 4193 1787 4207
rect 1853 4193 1867 4207
rect 1913 4193 1927 4207
rect 1953 4193 1967 4207
rect 1993 4193 2007 4207
rect 2053 4193 2067 4207
rect 2093 4193 2107 4207
rect 2493 4193 2507 4207
rect 2873 4193 2887 4207
rect 3013 4193 3027 4207
rect 3053 4193 3067 4207
rect 3113 4193 3127 4207
rect 3213 4193 3227 4207
rect 3293 4193 3307 4207
rect 3693 4193 3707 4207
rect 4173 4193 4187 4207
rect 4213 4193 4227 4207
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 153 4173 167 4187
rect 293 4173 307 4187
rect 333 4173 347 4187
rect 393 4173 407 4187
rect 433 4173 447 4187
rect 453 4173 467 4187
rect 493 4173 507 4187
rect 633 4173 647 4187
rect 893 4173 907 4187
rect 933 4173 947 4187
rect 973 4173 987 4187
rect 1573 4173 1587 4187
rect 1613 4173 1627 4187
rect 1653 4173 1667 4187
rect 1693 4173 1707 4187
rect 1713 4173 1727 4187
rect 1753 4173 1767 4187
rect 2233 4173 2247 4187
rect 2273 4173 2287 4187
rect 2353 4173 2367 4187
rect 2393 4173 2407 4187
rect 2433 4173 2447 4187
rect 2553 4173 2567 4187
rect 2593 4173 2607 4187
rect 2633 4173 2647 4187
rect 2713 4173 2727 4187
rect 2753 4173 2767 4187
rect 2933 4173 2947 4187
rect 2973 4173 2987 4187
rect 2993 4173 3007 4187
rect 3033 4173 3047 4187
rect 3333 4173 3347 4187
rect 3373 4173 3387 4187
rect 3493 4173 3507 4187
rect 3533 4173 3547 4187
rect 3613 4173 3627 4187
rect 3733 4173 3747 4187
rect 3773 4173 3787 4187
rect 3833 4173 3847 4187
rect 3913 4173 3927 4187
rect 3953 4173 3967 4187
rect 4053 4173 4067 4187
rect 4093 4173 4107 4187
rect 4153 4173 4167 4187
rect 4233 4173 4247 4187
rect 4273 4173 4287 4187
rect 4333 4173 4347 4187
rect 4373 4173 4387 4187
rect 4413 4173 4427 4187
rect 4513 4173 4527 4187
rect 4593 4173 4607 4187
rect 4633 4173 4647 4187
rect 113 4153 127 4167
rect 313 4153 327 4167
rect 593 4153 607 4167
rect 673 4153 687 4167
rect 753 4153 767 4167
rect 1593 4153 1607 4167
rect 1673 4153 1687 4167
rect 1893 4153 1907 4167
rect 2513 4153 2527 4167
rect 2573 4153 2587 4167
rect 2853 4153 2867 4167
rect 2953 4153 2967 4167
rect 3353 4153 3367 4167
rect 3753 4153 3767 4167
rect 4073 4153 4087 4167
rect 4193 4153 4207 4167
rect 4353 4153 4367 4167
rect 4453 4153 4467 4167
rect 373 4013 387 4027
rect 493 4013 507 4027
rect 1153 4013 1167 4027
rect 1273 4013 1287 4027
rect 1653 4013 1667 4027
rect 1913 4013 1927 4027
rect 2013 4013 2027 4027
rect 2133 4013 2147 4027
rect 2893 4013 2907 4027
rect 3073 4013 3087 4027
rect 3273 4013 3287 4027
rect 3453 4013 3467 4027
rect 3533 4013 3547 4027
rect 3853 4013 3867 4027
rect 3913 4013 3927 4027
rect 4013 4013 4027 4027
rect 4393 4013 4407 4027
rect 4653 4013 4667 4027
rect 293 3993 307 4007
rect 333 3993 347 4007
rect 413 3993 427 4007
rect 473 3993 487 4007
rect 513 3993 527 4007
rect 613 3993 627 4007
rect 653 3993 667 4007
rect 953 3993 967 4007
rect 993 3993 1007 4007
rect 1013 3993 1027 4007
rect 1053 3993 1067 4007
rect 1633 3993 1647 4007
rect 1673 3993 1687 4007
rect 1713 3993 1727 4007
rect 1773 3993 1787 4007
rect 1833 3993 1847 4007
rect 1873 3993 1887 4007
rect 1893 3993 1907 4007
rect 1933 3993 1947 4007
rect 2033 3993 2047 4007
rect 2073 3993 2087 4007
rect 2373 3993 2387 4007
rect 2413 3993 2427 4007
rect 2733 3993 2747 4007
rect 2773 3993 2787 4007
rect 2853 3993 2867 4007
rect 2953 3993 2967 4007
rect 2993 3993 3007 4007
rect 3053 3993 3067 4007
rect 3093 3993 3107 4007
rect 3233 3993 3247 4007
rect 3313 3993 3327 4007
rect 3373 3993 3387 4007
rect 3433 3993 3447 4007
rect 3473 3993 3487 4007
rect 3573 3993 3587 4007
rect 3653 3993 3667 4007
rect 3693 3993 3707 4007
rect 3813 3993 3827 4007
rect 3893 3993 3907 4007
rect 3933 3993 3947 4007
rect 3993 3993 4007 4007
rect 4033 3993 4047 4007
rect 4053 3993 4067 4007
rect 4113 3993 4127 4007
rect 4153 3993 4167 4007
rect 4193 3993 4207 4007
rect 4293 3993 4307 4007
rect 4333 3993 4347 4007
rect 4433 3993 4447 4007
rect 4513 3993 4527 4007
rect 4553 3993 4567 4007
rect 53 3973 67 3987
rect 113 3973 127 3987
rect 213 3973 227 3987
rect 273 3973 287 3987
rect 313 3973 327 3987
rect 353 3973 367 3987
rect 393 3973 407 3987
rect 553 3973 567 3987
rect 633 3973 647 3987
rect 673 3973 687 3987
rect 753 3973 767 3987
rect 793 3973 807 3987
rect 813 3973 827 3987
rect 853 3973 867 3987
rect 933 3973 947 3987
rect 973 3973 987 3987
rect 1033 3973 1047 3987
rect 1073 3973 1087 3987
rect 1133 3973 1147 3987
rect 1213 3973 1227 3987
rect 1253 3973 1267 3987
rect 1293 3973 1307 3987
rect 1333 3973 1347 3987
rect 1373 3973 1387 3987
rect 1433 3973 1447 3987
rect 1473 3973 1487 3987
rect 1553 3973 1567 3987
rect 1813 3973 1827 3987
rect 1853 3973 1867 3987
rect 1993 3973 2007 3987
rect 2053 3973 2067 3987
rect 2093 3973 2107 3987
rect 2153 3973 2167 3987
rect 2213 3973 2227 3987
rect 2273 3973 2287 3987
rect 2313 3973 2327 3987
rect 2473 3973 2487 3987
rect 2613 3973 2627 3987
rect 2913 3973 2927 3987
rect 2973 3973 2987 3987
rect 3013 3973 3027 3987
rect 3153 3973 3167 3987
rect 3253 3973 3267 3987
rect 3293 3973 3307 3987
rect 3513 3973 3527 3987
rect 3833 3973 3847 3987
rect 3873 3973 3887 3987
rect 4173 3973 4187 3987
rect 4213 3973 4227 3987
rect 4273 3973 4287 3987
rect 4313 3973 4327 3987
rect 4373 3973 4387 3987
rect 4673 3973 4687 3987
rect 33 3953 47 3967
rect 73 3953 87 3967
rect 93 3953 107 3967
rect 133 3953 147 3967
rect 193 3953 207 3967
rect 233 3953 247 3967
rect 533 3953 547 3967
rect 573 3953 587 3967
rect 733 3953 747 3967
rect 773 3953 787 3967
rect 833 3953 847 3967
rect 873 3953 887 3967
rect 1193 3953 1207 3967
rect 1233 3953 1247 3967
rect 1353 3953 1367 3967
rect 1393 3953 1407 3967
rect 1453 3953 1467 3967
rect 1493 3953 1507 3967
rect 1533 3953 1547 3967
rect 1573 3953 1587 3967
rect 1733 3953 1747 3967
rect 2193 3953 2207 3967
rect 2233 3953 2247 3967
rect 2293 3953 2307 3967
rect 2333 3953 2347 3967
rect 3133 3953 3147 3967
rect 3173 3953 3187 3967
rect 3353 3953 3367 3967
rect 4093 3953 4107 3967
rect 393 3733 407 3747
rect 473 3733 487 3747
rect 513 3733 527 3747
rect 553 3733 567 3747
rect 593 3733 607 3747
rect 773 3733 787 3747
rect 813 3733 827 3747
rect 873 3733 887 3747
rect 913 3733 927 3747
rect 1073 3733 1087 3747
rect 1113 3733 1127 3747
rect 1333 3733 1347 3747
rect 1373 3733 1387 3747
rect 1933 3733 1947 3747
rect 1973 3733 1987 3747
rect 3533 3733 3547 3747
rect 113 3713 127 3727
rect 153 3713 167 3727
rect 213 3713 227 3727
rect 293 3713 307 3727
rect 333 3713 347 3727
rect 493 3713 507 3727
rect 573 3713 587 3727
rect 633 3713 647 3727
rect 693 3713 707 3727
rect 733 3713 747 3727
rect 793 3713 807 3727
rect 893 3713 907 3727
rect 933 3713 947 3727
rect 953 3713 967 3727
rect 993 3713 1007 3727
rect 1053 3713 1067 3727
rect 1093 3713 1107 3727
rect 1153 3713 1167 3727
rect 1193 3713 1207 3727
rect 1273 3713 1287 3727
rect 1353 3713 1367 3727
rect 1393 3713 1407 3727
rect 1433 3713 1447 3727
rect 1493 3713 1507 3727
rect 1533 3713 1547 3727
rect 1593 3713 1607 3727
rect 1633 3713 1647 3727
rect 1673 3713 1687 3727
rect 1853 3713 1867 3727
rect 1893 3713 1907 3727
rect 1953 3713 1967 3727
rect 2053 3713 2067 3727
rect 2193 3713 2207 3727
rect 2333 3713 2347 3727
rect 2633 3713 2647 3727
rect 2673 3713 2687 3727
rect 2733 3713 2747 3727
rect 3033 3713 3047 3727
rect 3093 3713 3107 3727
rect 3153 3713 3167 3727
rect 3193 3713 3207 3727
rect 3273 3713 3287 3727
rect 3313 3713 3327 3727
rect 3333 3713 3347 3727
rect 3373 3713 3387 3727
rect 3453 3713 3467 3727
rect 3613 3713 3627 3727
rect 3653 3713 3667 3727
rect 3713 3713 3727 3727
rect 3753 3713 3767 3727
rect 4193 3713 4207 3727
rect 4233 3713 4247 3727
rect 4633 3713 4647 3727
rect 4693 3713 4707 3727
rect 33 3693 47 3707
rect 73 3693 87 3707
rect 93 3693 107 3707
rect 133 3693 147 3707
rect 273 3693 287 3707
rect 373 3693 387 3707
rect 433 3693 447 3707
rect 673 3693 687 3707
rect 713 3693 727 3707
rect 1013 3693 1027 3707
rect 1213 3693 1227 3707
rect 1513 3693 1527 3707
rect 1553 3693 1567 3707
rect 1693 3693 1707 3707
rect 1733 3693 1747 3707
rect 1773 3693 1787 3707
rect 1833 3693 1847 3707
rect 2013 3693 2027 3707
rect 2093 3693 2107 3707
rect 2133 3693 2147 3707
rect 2453 3693 2467 3707
rect 2493 3693 2507 3707
rect 2573 3693 2587 3707
rect 2653 3693 2667 3707
rect 2693 3693 2707 3707
rect 2793 3693 2807 3707
rect 2833 3693 2847 3707
rect 2873 3693 2887 3707
rect 2913 3693 2927 3707
rect 2953 3693 2967 3707
rect 2993 3693 3007 3707
rect 3133 3693 3147 3707
rect 3173 3693 3187 3707
rect 3253 3693 3267 3707
rect 3393 3693 3407 3707
rect 3493 3693 3507 3707
rect 3553 3693 3567 3707
rect 3593 3693 3607 3707
rect 3633 3693 3647 3707
rect 3693 3693 3707 3707
rect 3733 3693 3747 3707
rect 3873 3693 3887 3707
rect 3913 3693 3927 3707
rect 3993 3693 4007 3707
rect 4033 3693 4047 3707
rect 4073 3693 4087 3707
rect 4133 3693 4147 3707
rect 4173 3693 4187 3707
rect 4253 3693 4267 3707
rect 4313 3693 4327 3707
rect 4393 3693 4407 3707
rect 4433 3693 4447 3707
rect 4533 3693 4547 3707
rect 4573 3693 4587 3707
rect 53 3673 67 3687
rect 233 3673 247 3687
rect 313 3673 327 3687
rect 613 3673 627 3687
rect 973 3673 987 3687
rect 1173 3673 1187 3687
rect 1253 3673 1267 3687
rect 1453 3673 1467 3687
rect 1613 3673 1627 3687
rect 1653 3673 1667 3687
rect 1753 3673 1767 3687
rect 1873 3673 1887 3687
rect 1993 3673 2007 3687
rect 2753 3673 2767 3687
rect 2813 3673 2827 3687
rect 2893 3673 2907 3687
rect 2973 3673 2987 3687
rect 3013 3673 3027 3687
rect 3113 3673 3127 3687
rect 3293 3673 3307 3687
rect 3353 3673 3367 3687
rect 3433 3673 3447 3687
rect 4153 3673 4167 3687
rect 4213 3673 4227 3687
rect 4653 3673 4667 3687
rect 4673 3673 4687 3687
rect 373 3533 387 3547
rect 873 3533 887 3547
rect 1053 3533 1067 3547
rect 1153 3533 1167 3547
rect 2313 3533 2327 3547
rect 2373 3533 2387 3547
rect 3313 3533 3327 3547
rect 3353 3533 3367 3547
rect 3413 3533 3427 3547
rect 3513 3533 3527 3547
rect 3573 3533 3587 3547
rect 3653 3533 3667 3547
rect 173 3513 187 3527
rect 213 3513 227 3527
rect 293 3513 307 3527
rect 513 3513 527 3527
rect 553 3513 567 3527
rect 613 3513 627 3527
rect 653 3513 667 3527
rect 753 3513 767 3527
rect 793 3513 807 3527
rect 833 3513 847 3527
rect 1093 3513 1107 3527
rect 1133 3513 1147 3527
rect 1173 3513 1187 3527
rect 1373 3513 1387 3527
rect 1413 3513 1427 3527
rect 1553 3513 1567 3527
rect 1593 3513 1607 3527
rect 1673 3513 1687 3527
rect 1793 3513 1807 3527
rect 1833 3513 1847 3527
rect 1913 3513 1927 3527
rect 2053 3513 2067 3527
rect 2113 3513 2127 3527
rect 2453 3513 2467 3527
rect 2533 3513 2547 3527
rect 2573 3513 2587 3527
rect 2673 3513 2687 3527
rect 2713 3513 2727 3527
rect 2773 3513 2787 3527
rect 2813 3513 2827 3527
rect 2953 3513 2967 3527
rect 3033 3513 3047 3527
rect 3073 3513 3087 3527
rect 3213 3513 3227 3527
rect 3253 3513 3267 3527
rect 3333 3513 3347 3527
rect 3373 3513 3387 3527
rect 3493 3513 3507 3527
rect 3533 3513 3547 3527
rect 3613 3513 3627 3527
rect 3673 3513 3687 3527
rect 3773 3513 3787 3527
rect 3813 3513 3827 3527
rect 3853 3513 3867 3527
rect 3973 3513 3987 3527
rect 4053 3513 4067 3527
rect 4093 3513 4107 3527
rect 4213 3513 4227 3527
rect 4293 3513 4307 3527
rect 4333 3513 4347 3527
rect 4633 3513 4647 3527
rect 4673 3513 4687 3527
rect 53 3493 67 3507
rect 353 3493 367 3507
rect 433 3493 447 3507
rect 493 3493 507 3507
rect 533 3493 547 3507
rect 593 3493 607 3507
rect 633 3493 647 3507
rect 693 3493 707 3507
rect 773 3493 787 3507
rect 813 3493 827 3507
rect 893 3493 907 3507
rect 973 3493 987 3507
rect 1013 3493 1027 3507
rect 1033 3493 1047 3507
rect 1073 3493 1087 3507
rect 1233 3493 1247 3507
rect 1313 3493 1327 3507
rect 1393 3493 1407 3507
rect 1433 3493 1447 3507
rect 1753 3493 1767 3507
rect 1813 3493 1827 3507
rect 1853 3493 1867 3507
rect 1893 3493 1907 3507
rect 1993 3493 2007 3507
rect 2153 3493 2167 3507
rect 2213 3493 2227 3507
rect 2253 3493 2267 3507
rect 2333 3493 2347 3507
rect 2393 3493 2407 3507
rect 2693 3493 2707 3507
rect 2733 3493 2747 3507
rect 2873 3493 2887 3507
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3293 3493 3307 3507
rect 3433 3493 3447 3507
rect 3553 3493 3567 3507
rect 3593 3493 3607 3507
rect 3713 3493 3727 3507
rect 3793 3493 3807 3507
rect 3833 3493 3847 3507
rect 3913 3493 3927 3507
rect 4453 3493 4467 3507
rect 4593 3493 4607 3507
rect 4653 3493 4667 3507
rect 4693 3493 4707 3507
rect 33 3473 47 3487
rect 73 3473 87 3487
rect 413 3473 427 3487
rect 453 3473 467 3487
rect 673 3473 687 3487
rect 713 3473 727 3487
rect 953 3473 967 3487
rect 993 3473 1007 3487
rect 1213 3473 1227 3487
rect 1253 3473 1267 3487
rect 1293 3473 1307 3487
rect 1333 3473 1347 3487
rect 1733 3473 1747 3487
rect 1773 3473 1787 3487
rect 1973 3473 1987 3487
rect 2013 3473 2027 3487
rect 2073 3473 2087 3487
rect 2133 3473 2147 3487
rect 2173 3473 2187 3487
rect 2233 3473 2247 3487
rect 2273 3473 2287 3487
rect 2853 3473 2867 3487
rect 2893 3473 2907 3487
rect 3893 3473 3907 3487
rect 3933 3473 3947 3487
rect 393 3253 407 3267
rect 433 3253 447 3267
rect 913 3253 927 3267
rect 953 3253 967 3267
rect 1013 3253 1027 3267
rect 1053 3253 1067 3267
rect 1133 3253 1147 3267
rect 1213 3253 1227 3267
rect 1253 3253 1267 3267
rect 1393 3253 1407 3267
rect 1433 3253 1447 3267
rect 1593 3253 1607 3267
rect 1633 3253 1647 3267
rect 1853 3253 1867 3267
rect 1893 3253 1907 3267
rect 2353 3253 2367 3267
rect 2393 3253 2407 3267
rect 3493 3253 3507 3267
rect 3533 3253 3547 3267
rect 3573 3253 3587 3267
rect 3613 3253 3627 3267
rect 3653 3253 3667 3267
rect 3693 3253 3707 3267
rect 3733 3253 3747 3267
rect 3773 3253 3787 3267
rect 3913 3253 3927 3267
rect 3953 3253 3967 3267
rect 4473 3253 4487 3267
rect 4513 3253 4527 3267
rect 293 3233 307 3247
rect 333 3233 347 3247
rect 413 3233 427 3247
rect 713 3233 727 3247
rect 753 3233 767 3247
rect 833 3233 847 3247
rect 873 3233 887 3247
rect 933 3233 947 3247
rect 1033 3233 1047 3247
rect 1073 3233 1087 3247
rect 1193 3233 1207 3247
rect 1233 3233 1247 3247
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1413 3233 1427 3247
rect 1493 3233 1507 3247
rect 1613 3233 1627 3247
rect 1673 3233 1687 3247
rect 1713 3233 1727 3247
rect 1773 3233 1787 3247
rect 1813 3233 1827 3247
rect 1873 3233 1887 3247
rect 1953 3233 1967 3247
rect 1993 3233 2007 3247
rect 2053 3233 2067 3247
rect 2093 3233 2107 3247
rect 2153 3233 2167 3247
rect 2213 3233 2227 3247
rect 2253 3233 2267 3247
rect 2313 3233 2327 3247
rect 2373 3233 2387 3247
rect 3013 3233 3027 3247
rect 3053 3233 3067 3247
rect 3113 3233 3127 3247
rect 3153 3233 3167 3247
rect 3213 3233 3227 3247
rect 3253 3233 3267 3247
rect 3313 3233 3327 3247
rect 3353 3233 3367 3247
rect 3413 3233 3427 3247
rect 3453 3233 3467 3247
rect 3513 3233 3527 3247
rect 3593 3233 3607 3247
rect 3673 3233 3687 3247
rect 3753 3233 3767 3247
rect 3933 3233 3947 3247
rect 4153 3233 4167 3247
rect 4213 3233 4227 3247
rect 4253 3233 4267 3247
rect 4313 3233 4327 3247
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4493 3233 4507 3247
rect 93 3213 107 3227
rect 133 3213 147 3227
rect 213 3213 227 3227
rect 273 3213 287 3227
rect 313 3213 327 3227
rect 353 3213 367 3227
rect 473 3213 487 3227
rect 553 3213 567 3227
rect 593 3213 607 3227
rect 733 3213 747 3227
rect 773 3213 787 3227
rect 813 3213 827 3227
rect 853 3213 867 3227
rect 893 3213 907 3227
rect 1113 3213 1127 3227
rect 1173 3213 1187 3227
rect 1293 3213 1307 3227
rect 1333 3213 1347 3227
rect 1533 3213 1547 3227
rect 1653 3213 1667 3227
rect 1693 3213 1707 3227
rect 1793 3213 1807 3227
rect 1833 3213 1847 3227
rect 1933 3213 1947 3227
rect 1973 3213 1987 3227
rect 2073 3213 2087 3227
rect 2113 3213 2127 3227
rect 2193 3213 2207 3227
rect 2233 3213 2247 3227
rect 2453 3213 2467 3227
rect 2533 3213 2547 3227
rect 2573 3213 2587 3227
rect 2673 3213 2687 3227
rect 2713 3213 2727 3227
rect 2773 3213 2787 3227
rect 2853 3213 2867 3227
rect 2893 3213 2907 3227
rect 3033 3213 3047 3227
rect 3073 3213 3087 3227
rect 3133 3213 3147 3227
rect 3173 3213 3187 3227
rect 3193 3213 3207 3227
rect 3233 3213 3247 3227
rect 3333 3213 3347 3227
rect 3373 3213 3387 3227
rect 3393 3213 3407 3227
rect 3433 3213 3447 3227
rect 3813 3213 3827 3227
rect 3853 3213 3867 3227
rect 3993 3213 4007 3227
rect 4033 3213 4047 3227
rect 4053 3213 4067 3227
rect 4093 3213 4107 3227
rect 4233 3213 4247 3227
rect 4273 3213 4287 3227
rect 4353 3213 4367 3227
rect 4393 3213 4407 3227
rect 4613 3213 4627 3227
rect 4653 3213 4667 3227
rect 4733 3213 4747 3227
rect 1553 3193 1567 3207
rect 2133 3193 2147 3207
rect 2333 3193 2347 3207
rect 4013 3193 4027 3207
rect 4173 3193 4187 3207
rect 4333 3193 4347 3207
rect 773 3053 787 3067
rect 1133 3053 1147 3067
rect 1873 3053 1887 3067
rect 1953 3053 1967 3067
rect 2033 3053 2047 3067
rect 2213 3053 2227 3067
rect 2453 3053 2467 3067
rect 3053 3053 3067 3067
rect 3153 3053 3167 3067
rect 3213 3053 3227 3067
rect 3773 3053 3787 3067
rect 4233 3053 4247 3067
rect 33 3033 47 3047
rect 73 3033 87 3047
rect 113 3033 127 3047
rect 153 3033 167 3047
rect 213 3033 227 3047
rect 253 3033 267 3047
rect 333 3033 347 3047
rect 373 3033 387 3047
rect 473 3033 487 3047
rect 513 3033 527 3047
rect 753 3033 767 3047
rect 793 3033 807 3047
rect 933 3033 947 3047
rect 973 3033 987 3047
rect 1033 3033 1047 3047
rect 1073 3033 1087 3047
rect 1113 3033 1127 3047
rect 1153 3033 1167 3047
rect 1213 3033 1227 3047
rect 1253 3033 1267 3047
rect 1373 3033 1387 3047
rect 1573 3033 1587 3047
rect 1613 3033 1627 3047
rect 1653 3033 1667 3047
rect 1693 3033 1707 3047
rect 1753 3033 1767 3047
rect 1793 3033 1807 3047
rect 1853 3033 1867 3047
rect 1893 3033 1907 3047
rect 1993 3033 2007 3047
rect 2093 3033 2107 3047
rect 2133 3033 2147 3047
rect 2193 3033 2207 3047
rect 2233 3033 2247 3047
rect 2353 3033 2367 3047
rect 2393 3033 2407 3047
rect 2513 3033 2527 3047
rect 2553 3033 2567 3047
rect 2613 3033 2627 3047
rect 2653 3033 2667 3047
rect 2853 3033 2867 3047
rect 2893 3033 2907 3047
rect 2973 3033 2987 3047
rect 3033 3033 3047 3047
rect 3073 3033 3087 3047
rect 3113 3033 3127 3047
rect 3193 3033 3207 3047
rect 3233 3033 3247 3047
rect 3353 3033 3367 3047
rect 3393 3033 3407 3047
rect 3473 3033 3487 3047
rect 3593 3033 3607 3047
rect 3633 3033 3647 3047
rect 3713 3033 3727 3047
rect 3753 3033 3767 3047
rect 3793 3033 3807 3047
rect 3873 3033 3887 3047
rect 3913 3033 3927 3047
rect 3973 3033 3987 3047
rect 4013 3033 4027 3047
rect 4033 3033 4047 3047
rect 4073 3033 4087 3047
rect 4133 3033 4147 3047
rect 4173 3033 4187 3047
rect 4413 3033 4427 3047
rect 4493 3033 4507 3047
rect 4533 3033 4547 3047
rect 4633 3033 4647 3047
rect 4673 3033 4687 3047
rect 53 3013 67 3027
rect 93 3013 107 3027
rect 493 3013 507 3027
rect 533 3013 547 3027
rect 593 3013 607 3027
rect 693 3013 707 3027
rect 833 3013 847 3027
rect 913 3013 927 3027
rect 953 3013 967 3027
rect 1013 3013 1027 3027
rect 1053 3013 1067 3027
rect 1193 3013 1207 3027
rect 1233 3013 1247 3027
rect 1293 3013 1307 3027
rect 1393 3013 1407 3027
rect 1433 3013 1447 3027
rect 1513 3013 1527 3027
rect 1673 3013 1687 3027
rect 1713 3013 1727 3027
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1933 3013 1947 3027
rect 1973 3013 1987 3027
rect 2053 3013 2067 3027
rect 2113 3013 2127 3027
rect 2153 3013 2167 3027
rect 2313 3013 2327 3027
rect 2373 3013 2387 3027
rect 2413 3013 2427 3027
rect 2473 3013 2487 3027
rect 2533 3013 2547 3027
rect 2573 3013 2587 3027
rect 2713 3013 2727 3027
rect 3133 3013 3147 3027
rect 3173 3013 3187 3027
rect 3853 3013 3867 3027
rect 3893 3013 3907 3027
rect 3953 3013 3967 3027
rect 3993 3013 4007 3027
rect 4053 3013 4067 3027
rect 4093 3013 4107 3027
rect 4153 3013 4167 3027
rect 4193 3013 4207 3027
rect 4253 3013 4267 3027
rect 4293 3013 4307 3027
rect 4333 3013 4347 3027
rect 4653 3013 4667 3027
rect 4693 3013 4707 3027
rect 173 2993 187 3007
rect 573 2993 587 3007
rect 613 2993 627 3007
rect 673 2993 687 3007
rect 713 2993 727 3007
rect 813 2993 827 3007
rect 853 2993 867 3007
rect 1273 2993 1287 3007
rect 1313 2993 1327 3007
rect 1413 2993 1427 3007
rect 1453 2993 1467 3007
rect 1493 2993 1507 3007
rect 1533 2993 1547 3007
rect 2293 2993 2307 3007
rect 2333 2993 2347 3007
rect 2693 2993 2707 3007
rect 2733 2993 2747 3007
rect 4313 2993 4327 3007
rect 4353 2993 4367 3007
rect 293 2773 307 2787
rect 333 2773 347 2787
rect 413 2773 427 2787
rect 573 2773 587 2787
rect 613 2773 627 2787
rect 773 2773 787 2787
rect 813 2773 827 2787
rect 893 2773 907 2787
rect 1053 2773 1067 2787
rect 1093 2773 1107 2787
rect 2553 2773 2567 2787
rect 2813 2773 2827 2787
rect 2853 2773 2867 2787
rect 4633 2773 4647 2787
rect 4673 2773 4687 2787
rect 33 2753 47 2767
rect 93 2753 107 2767
rect 133 2753 147 2767
rect 193 2753 207 2767
rect 233 2753 247 2767
rect 313 2753 327 2767
rect 493 2753 507 2767
rect 533 2753 547 2767
rect 593 2753 607 2767
rect 693 2753 707 2767
rect 753 2753 767 2767
rect 793 2753 807 2767
rect 973 2753 987 2767
rect 1013 2753 1027 2767
rect 1073 2753 1087 2767
rect 1153 2753 1167 2767
rect 1193 2753 1207 2767
rect 1813 2753 1827 2767
rect 1853 2753 1867 2767
rect 1913 2753 1927 2767
rect 1973 2753 1987 2767
rect 2013 2753 2027 2767
rect 2333 2753 2347 2767
rect 2473 2753 2487 2767
rect 2633 2753 2647 2767
rect 2673 2753 2687 2767
rect 2733 2753 2747 2767
rect 2773 2753 2787 2767
rect 2833 2753 2847 2767
rect 3393 2753 3407 2767
rect 3553 2753 3567 2767
rect 3853 2753 3867 2767
rect 3893 2753 3907 2767
rect 4033 2753 4047 2767
rect 4073 2753 4087 2767
rect 4133 2753 4147 2767
rect 4173 2753 4187 2767
rect 4553 2753 4567 2767
rect 4593 2753 4607 2767
rect 4653 2753 4667 2767
rect 113 2733 127 2747
rect 153 2733 167 2747
rect 173 2733 187 2747
rect 213 2733 227 2747
rect 253 2733 267 2747
rect 373 2733 387 2747
rect 433 2733 447 2747
rect 513 2733 527 2747
rect 553 2733 567 2747
rect 673 2733 687 2747
rect 733 2733 747 2747
rect 853 2733 867 2747
rect 913 2733 927 2747
rect 993 2733 1007 2747
rect 1033 2733 1047 2747
rect 1173 2733 1187 2747
rect 1213 2733 1227 2747
rect 1253 2733 1267 2747
rect 1333 2733 1347 2747
rect 1373 2733 1387 2747
rect 1493 2733 1507 2747
rect 1533 2733 1547 2747
rect 1633 2733 1647 2747
rect 1673 2733 1687 2747
rect 1753 2733 1767 2747
rect 1793 2733 1807 2747
rect 1833 2733 1847 2747
rect 1953 2733 1967 2747
rect 1993 2733 2007 2747
rect 2033 2733 2047 2747
rect 2093 2733 2107 2747
rect 2133 2733 2147 2747
rect 2173 2733 2187 2747
rect 2213 2733 2227 2747
rect 2253 2733 2267 2747
rect 2293 2733 2307 2747
rect 2393 2733 2407 2747
rect 2433 2733 2447 2747
rect 2513 2733 2527 2747
rect 2573 2733 2587 2747
rect 2613 2733 2627 2747
rect 2653 2733 2667 2747
rect 2713 2733 2727 2747
rect 2753 2733 2767 2747
rect 2973 2733 2987 2747
rect 3013 2733 3027 2747
rect 3093 2733 3107 2747
rect 3213 2733 3227 2747
rect 3253 2733 3267 2747
rect 3333 2733 3347 2747
rect 3453 2733 3467 2747
rect 3493 2733 3507 2747
rect 3533 2733 3547 2747
rect 3653 2733 3667 2747
rect 3693 2733 3707 2747
rect 3773 2733 3787 2747
rect 3833 2733 3847 2747
rect 3873 2733 3887 2747
rect 3913 2733 3927 2747
rect 3953 2733 3967 2747
rect 3993 2733 4007 2747
rect 4013 2733 4027 2747
rect 4053 2733 4067 2747
rect 4153 2733 4167 2747
rect 4193 2733 4207 2747
rect 4213 2733 4227 2747
rect 4253 2733 4267 2747
rect 4373 2733 4387 2747
rect 4413 2733 4427 2747
rect 4493 2733 4507 2747
rect 4533 2733 4547 2747
rect 4573 2733 4587 2747
rect 53 2713 67 2727
rect 1893 2713 1907 2727
rect 2113 2713 2127 2727
rect 2193 2713 2207 2727
rect 2273 2713 2287 2727
rect 2313 2713 2327 2727
rect 2413 2713 2427 2727
rect 2453 2713 2467 2727
rect 3413 2713 3427 2727
rect 3473 2713 3487 2727
rect 3973 2713 3987 2727
rect 4233 2713 4247 2727
rect 133 2573 147 2587
rect 253 2573 267 2587
rect 433 2573 447 2587
rect 1233 2573 1247 2587
rect 2093 2573 2107 2587
rect 2193 2573 2207 2587
rect 2253 2573 2267 2587
rect 2333 2573 2347 2587
rect 2473 2573 2487 2587
rect 2813 2573 2827 2587
rect 3913 2573 3927 2587
rect 3973 2573 3987 2587
rect 173 2553 187 2567
rect 293 2553 307 2567
rect 353 2553 367 2567
rect 393 2553 407 2567
rect 613 2553 627 2567
rect 653 2553 667 2567
rect 693 2553 707 2567
rect 953 2553 967 2567
rect 993 2553 1007 2567
rect 1293 2553 1307 2567
rect 1333 2553 1347 2567
rect 1453 2553 1467 2567
rect 1653 2553 1667 2567
rect 1693 2553 1707 2567
rect 1773 2553 1787 2567
rect 2073 2553 2087 2567
rect 2113 2553 2127 2567
rect 2233 2553 2247 2567
rect 2273 2553 2287 2567
rect 2393 2553 2407 2567
rect 2433 2553 2447 2567
rect 2453 2553 2467 2567
rect 2493 2553 2507 2567
rect 2533 2553 2547 2567
rect 2593 2553 2607 2567
rect 2633 2553 2647 2567
rect 2673 2553 2687 2567
rect 2833 2553 2847 2567
rect 2993 2553 3007 2567
rect 3033 2553 3047 2567
rect 3073 2553 3087 2567
rect 3113 2553 3127 2567
rect 3193 2553 3207 2567
rect 3233 2553 3247 2567
rect 3333 2553 3347 2567
rect 3373 2553 3387 2567
rect 3413 2553 3427 2567
rect 3453 2553 3467 2567
rect 3493 2553 3507 2567
rect 3553 2553 3567 2567
rect 3593 2553 3607 2567
rect 3693 2553 3707 2567
rect 3733 2553 3747 2567
rect 3813 2553 3827 2567
rect 3873 2553 3887 2567
rect 3953 2553 3967 2567
rect 3993 2553 4007 2567
rect 4313 2553 4327 2567
rect 4353 2553 4367 2567
rect 4433 2553 4447 2567
rect 4473 2553 4487 2567
rect 4513 2553 4527 2567
rect 13 2533 27 2547
rect 53 2533 67 2547
rect 113 2533 127 2547
rect 153 2533 167 2547
rect 233 2533 247 2547
rect 413 2533 427 2547
rect 453 2533 467 2547
rect 513 2533 527 2547
rect 553 2533 567 2547
rect 593 2533 607 2547
rect 633 2533 647 2547
rect 713 2533 727 2547
rect 773 2533 787 2547
rect 853 2533 867 2547
rect 893 2533 907 2547
rect 933 2533 947 2547
rect 973 2533 987 2547
rect 1033 2533 1047 2547
rect 1133 2533 1147 2547
rect 1173 2533 1187 2547
rect 1213 2533 1227 2547
rect 1273 2533 1287 2547
rect 1313 2533 1327 2547
rect 1373 2533 1387 2547
rect 1433 2533 1447 2547
rect 1533 2533 1547 2547
rect 1833 2533 1847 2547
rect 1913 2533 1927 2547
rect 1973 2533 1987 2547
rect 2013 2533 2027 2547
rect 2173 2533 2187 2547
rect 2313 2533 2327 2547
rect 2373 2533 2387 2547
rect 2413 2533 2427 2547
rect 2653 2533 2667 2547
rect 2693 2533 2707 2547
rect 2773 2533 2787 2547
rect 2873 2533 2887 2547
rect 2933 2533 2947 2547
rect 3093 2533 3107 2547
rect 3133 2533 3147 2547
rect 3293 2533 3307 2547
rect 3353 2533 3367 2547
rect 3393 2533 3407 2547
rect 3893 2533 3907 2547
rect 3933 2533 3947 2547
rect 4053 2533 4067 2547
rect 4193 2533 4207 2547
rect 4493 2533 4507 2547
rect 4533 2533 4547 2547
rect 4593 2533 4607 2547
rect 4673 2533 4687 2547
rect 33 2513 47 2527
rect 73 2513 87 2527
rect 313 2513 327 2527
rect 493 2513 507 2527
rect 533 2513 547 2527
rect 753 2513 767 2527
rect 793 2513 807 2527
rect 833 2513 847 2527
rect 873 2513 887 2527
rect 1013 2513 1027 2527
rect 1053 2513 1067 2527
rect 1113 2513 1127 2527
rect 1153 2513 1167 2527
rect 1353 2513 1367 2527
rect 1393 2513 1407 2527
rect 1513 2513 1527 2527
rect 1553 2513 1567 2527
rect 1813 2513 1827 2527
rect 1853 2513 1867 2527
rect 1893 2513 1907 2527
rect 1933 2513 1947 2527
rect 1993 2513 2007 2527
rect 2033 2513 2047 2527
rect 2573 2513 2587 2527
rect 2753 2513 2767 2527
rect 2793 2513 2807 2527
rect 2913 2513 2927 2527
rect 2953 2513 2967 2527
rect 3273 2513 3287 2527
rect 3313 2513 3327 2527
rect 4573 2513 4587 2527
rect 4613 2513 4627 2527
rect 4653 2513 4667 2527
rect 4693 2513 4707 2527
rect 33 2293 47 2307
rect 73 2293 87 2307
rect 333 2293 347 2307
rect 373 2293 387 2307
rect 813 2293 827 2307
rect 873 2293 887 2307
rect 913 2293 927 2307
rect 993 2293 1007 2307
rect 2513 2293 2527 2307
rect 2553 2293 2567 2307
rect 2633 2293 2647 2307
rect 3773 2293 3787 2307
rect 3813 2293 3827 2307
rect 4653 2293 4667 2307
rect 4693 2293 4707 2307
rect 53 2273 67 2287
rect 93 2273 107 2287
rect 133 2273 147 2287
rect 173 2273 187 2287
rect 233 2273 247 2287
rect 273 2273 287 2287
rect 313 2273 327 2287
rect 353 2273 367 2287
rect 413 2273 427 2287
rect 453 2273 467 2287
rect 533 2273 547 2287
rect 573 2273 587 2287
rect 653 2273 667 2287
rect 693 2273 707 2287
rect 733 2273 747 2287
rect 893 2273 907 2287
rect 1073 2273 1087 2287
rect 1113 2273 1127 2287
rect 1173 2273 1187 2287
rect 1213 2273 1227 2287
rect 1513 2273 1527 2287
rect 1553 2273 1567 2287
rect 1853 2273 1867 2287
rect 1913 2273 1927 2287
rect 1973 2273 1987 2287
rect 2013 2273 2027 2287
rect 2333 2273 2347 2287
rect 2373 2273 2387 2287
rect 2433 2273 2447 2287
rect 2473 2273 2487 2287
rect 2493 2273 2507 2287
rect 2533 2273 2547 2287
rect 2953 2273 2967 2287
rect 2993 2273 3007 2287
rect 3053 2273 3067 2287
rect 3093 2273 3107 2287
rect 3153 2273 3167 2287
rect 3193 2273 3207 2287
rect 3493 2273 3507 2287
rect 3533 2273 3547 2287
rect 3713 2273 3727 2287
rect 3793 2273 3807 2287
rect 3873 2273 3887 2287
rect 3913 2273 3927 2287
rect 3993 2273 4007 2287
rect 4033 2273 4047 2287
rect 4573 2273 4587 2287
rect 4613 2273 4627 2287
rect 4673 2273 4687 2287
rect 153 2253 167 2267
rect 193 2253 207 2267
rect 213 2253 227 2267
rect 253 2253 267 2267
rect 473 2253 487 2267
rect 513 2253 527 2267
rect 553 2253 567 2267
rect 633 2253 647 2267
rect 793 2253 807 2267
rect 853 2253 867 2267
rect 953 2253 967 2267
rect 1013 2253 1027 2267
rect 1093 2253 1107 2267
rect 1133 2253 1147 2267
rect 1193 2253 1207 2267
rect 1233 2253 1247 2267
rect 1333 2253 1347 2267
rect 1373 2253 1387 2267
rect 1453 2253 1467 2267
rect 1533 2253 1547 2267
rect 1573 2253 1587 2267
rect 1673 2253 1687 2267
rect 1713 2253 1727 2267
rect 1793 2253 1807 2267
rect 1953 2253 1967 2267
rect 1993 2253 2007 2267
rect 2133 2253 2147 2267
rect 2173 2253 2187 2267
rect 2253 2253 2267 2267
rect 2313 2253 2327 2267
rect 2413 2253 2427 2267
rect 2593 2253 2607 2267
rect 2653 2253 2667 2267
rect 2713 2253 2727 2267
rect 2793 2253 2807 2267
rect 2833 2253 2847 2267
rect 2973 2253 2987 2267
rect 3013 2253 3027 2267
rect 3073 2253 3087 2267
rect 3113 2253 3127 2267
rect 3133 2253 3147 2267
rect 3173 2253 3187 2267
rect 3253 2253 3267 2267
rect 3333 2253 3347 2267
rect 3373 2253 3387 2267
rect 3513 2253 3527 2267
rect 3553 2253 3567 2267
rect 3593 2253 3607 2267
rect 3633 2253 3647 2267
rect 3673 2253 3687 2267
rect 3853 2253 3867 2267
rect 3893 2253 3907 2267
rect 3933 2253 3947 2267
rect 3973 2253 3987 2267
rect 4013 2253 4027 2267
rect 4053 2253 4067 2267
rect 4153 2253 4167 2267
rect 4193 2253 4207 2267
rect 4273 2253 4287 2267
rect 4333 2253 4347 2267
rect 4413 2253 4427 2267
rect 4453 2253 4467 2267
rect 4553 2253 4567 2267
rect 4593 2253 4607 2267
rect 433 2233 447 2247
rect 673 2233 687 2247
rect 713 2233 727 2247
rect 1873 2233 1887 2247
rect 1933 2233 1947 2247
rect 2353 2233 2367 2247
rect 2453 2233 2467 2247
rect 3613 2233 3627 2247
rect 3653 2233 3667 2247
rect 313 2093 327 2107
rect 413 2093 427 2107
rect 713 2093 727 2107
rect 1213 2093 1227 2107
rect 1313 2093 1327 2107
rect 1733 2093 1747 2107
rect 1833 2093 1847 2107
rect 2573 2093 2587 2107
rect 3133 2093 3147 2107
rect 3193 2093 3207 2107
rect 4313 2093 4327 2107
rect 4413 2093 4427 2107
rect 4493 2093 4507 2107
rect 33 2073 47 2087
rect 73 2073 87 2087
rect 133 2073 147 2087
rect 173 2073 187 2087
rect 353 2073 367 2087
rect 453 2073 467 2087
rect 753 2073 767 2087
rect 833 2073 847 2087
rect 873 2073 887 2087
rect 1253 2073 1267 2087
rect 1293 2073 1307 2087
rect 1333 2073 1347 2087
rect 1653 2073 1667 2087
rect 1693 2073 1707 2087
rect 1773 2073 1787 2087
rect 1813 2073 1827 2087
rect 1853 2073 1867 2087
rect 1933 2073 1947 2087
rect 1973 2073 1987 2087
rect 1993 2073 2007 2087
rect 2033 2073 2047 2087
rect 2133 2073 2147 2087
rect 2173 2073 2187 2087
rect 2493 2073 2507 2087
rect 2553 2073 2567 2087
rect 2593 2073 2607 2087
rect 2913 2073 2927 2087
rect 2953 2073 2967 2087
rect 3033 2073 3047 2087
rect 3093 2073 3107 2087
rect 3173 2073 3187 2087
rect 3213 2073 3227 2087
rect 3273 2073 3287 2087
rect 3313 2073 3327 2087
rect 3353 2073 3367 2087
rect 3453 2073 3467 2087
rect 3493 2073 3507 2087
rect 3573 2073 3587 2087
rect 3613 2073 3627 2087
rect 3653 2073 3667 2087
rect 3793 2073 3807 2087
rect 3833 2073 3847 2087
rect 3913 2073 3927 2087
rect 3973 2073 3987 2087
rect 4053 2073 4067 2087
rect 4093 2073 4107 2087
rect 4213 2073 4227 2087
rect 4253 2073 4267 2087
rect 4293 2073 4307 2087
rect 4393 2073 4407 2087
rect 4433 2073 4447 2087
rect 4473 2073 4487 2087
rect 4513 2073 4527 2087
rect 4553 2073 4567 2087
rect 4633 2073 4647 2087
rect 4673 2073 4687 2087
rect 113 2053 127 2067
rect 153 2053 167 2067
rect 233 2053 247 2067
rect 273 2053 287 2067
rect 293 2053 307 2067
rect 333 2053 347 2067
rect 393 2053 407 2067
rect 433 2053 447 2067
rect 493 2053 507 2067
rect 533 2053 547 2067
rect 593 2053 607 2067
rect 633 2053 647 2067
rect 693 2053 707 2067
rect 733 2053 747 2067
rect 813 2053 827 2067
rect 853 2053 867 2067
rect 893 2053 907 2067
rect 933 2053 947 2067
rect 993 2053 1007 2067
rect 1033 2053 1047 2067
rect 1093 2053 1107 2067
rect 1133 2053 1147 2067
rect 1193 2053 1207 2067
rect 1233 2053 1247 2067
rect 1413 2053 1427 2067
rect 1493 2053 1507 2067
rect 1553 2053 1567 2067
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1713 2053 1727 2067
rect 1753 2053 1767 2067
rect 1913 2053 1927 2067
rect 1953 2053 1967 2067
rect 2013 2053 2027 2067
rect 2053 2053 2067 2067
rect 2113 2053 2127 2067
rect 2153 2053 2167 2067
rect 2213 2053 2227 2067
rect 2353 2053 2367 2067
rect 2413 2053 2427 2067
rect 2633 2053 2647 2067
rect 2713 2053 2727 2067
rect 2773 2053 2787 2067
rect 3113 2053 3127 2067
rect 3153 2053 3167 2067
rect 3293 2053 3307 2067
rect 3333 2053 3347 2067
rect 3633 2053 3647 2067
rect 3673 2053 3687 2067
rect 4233 2053 4247 2067
rect 4273 2053 4287 2067
rect 4333 2053 4347 2067
rect 213 2033 227 2047
rect 253 2033 267 2047
rect 513 2033 527 2047
rect 553 2033 567 2047
rect 613 2033 627 2047
rect 653 2033 667 2047
rect 913 2033 927 2047
rect 953 2033 967 2047
rect 1013 2033 1027 2047
rect 1053 2033 1067 2047
rect 1113 2033 1127 2047
rect 1153 2033 1167 2047
rect 1393 2033 1407 2047
rect 1433 2033 1447 2047
rect 1473 2033 1487 2047
rect 1513 2033 1527 2047
rect 1533 2033 1547 2047
rect 1573 2033 1587 2047
rect 2393 2033 2407 2047
rect 2433 2033 2447 2047
rect 2513 2033 2527 2047
rect 2693 2033 2707 2047
rect 2733 2033 2747 2047
rect 2753 2033 2767 2047
rect 2793 2033 2807 2047
rect 233 1813 247 1827
rect 273 1813 287 1827
rect 333 1813 347 1827
rect 373 1813 387 1827
rect 573 1813 587 1827
rect 993 1813 1007 1827
rect 1033 1813 1047 1827
rect 1153 1813 1167 1827
rect 1193 1813 1207 1827
rect 1253 1813 1267 1827
rect 1293 1813 1307 1827
rect 1533 1813 1547 1827
rect 1573 1813 1587 1827
rect 1753 1813 1767 1827
rect 1793 1813 1807 1827
rect 1873 1813 1887 1827
rect 2693 1813 2707 1827
rect 2733 1813 2747 1827
rect 3413 1813 3427 1827
rect 3453 1813 3467 1827
rect 3833 1813 3847 1827
rect 3873 1813 3887 1827
rect 4693 1813 4707 1827
rect 4733 1813 4747 1827
rect 53 1793 67 1807
rect 93 1793 107 1807
rect 153 1793 167 1807
rect 193 1793 207 1807
rect 253 1793 267 1807
rect 353 1793 367 1807
rect 393 1793 407 1807
rect 433 1793 447 1807
rect 473 1793 487 1807
rect 673 1793 687 1807
rect 793 1793 807 1807
rect 833 1793 847 1807
rect 893 1793 907 1807
rect 933 1793 947 1807
rect 973 1793 987 1807
rect 1013 1793 1027 1807
rect 1093 1793 1107 1807
rect 1133 1793 1147 1807
rect 1173 1793 1187 1807
rect 1233 1793 1247 1807
rect 1273 1793 1287 1807
rect 1353 1793 1367 1807
rect 1433 1793 1447 1807
rect 1473 1793 1487 1807
rect 1513 1793 1527 1807
rect 1553 1793 1567 1807
rect 1633 1793 1647 1807
rect 1713 1793 1727 1807
rect 1773 1793 1787 1807
rect 1813 1793 1827 1807
rect 2273 1793 2287 1807
rect 2333 1793 2347 1807
rect 2373 1793 2387 1807
rect 2593 1793 2607 1807
rect 2633 1793 2647 1807
rect 2713 1793 2727 1807
rect 2853 1793 2867 1807
rect 2893 1793 2907 1807
rect 2953 1793 2967 1807
rect 3333 1793 3347 1807
rect 3373 1793 3387 1807
rect 3433 1793 3447 1807
rect 3853 1793 3867 1807
rect 3913 1793 3927 1807
rect 3953 1793 3967 1807
rect 4013 1793 4027 1807
rect 4053 1793 4067 1807
rect 4153 1793 4167 1807
rect 4213 1793 4227 1807
rect 4253 1793 4267 1807
rect 4293 1793 4307 1807
rect 4713 1793 4727 1807
rect 33 1773 47 1787
rect 73 1773 87 1787
rect 113 1773 127 1787
rect 133 1773 147 1787
rect 173 1773 187 1787
rect 413 1773 427 1787
rect 453 1773 467 1787
rect 493 1773 507 1787
rect 533 1773 547 1787
rect 593 1773 607 1787
rect 653 1773 667 1787
rect 693 1773 707 1787
rect 733 1773 747 1787
rect 813 1773 827 1787
rect 853 1773 867 1787
rect 873 1773 887 1787
rect 913 1773 927 1787
rect 1413 1773 1427 1787
rect 1453 1773 1467 1787
rect 1493 1773 1507 1787
rect 1693 1773 1707 1787
rect 1833 1773 1847 1787
rect 1893 1773 1907 1787
rect 2013 1773 2027 1787
rect 2053 1773 2067 1787
rect 2133 1773 2147 1787
rect 2193 1773 2207 1787
rect 2233 1773 2247 1787
rect 2313 1773 2327 1787
rect 2353 1773 2367 1787
rect 2413 1773 2427 1787
rect 2453 1773 2467 1787
rect 2493 1773 2507 1787
rect 2533 1773 2547 1787
rect 2573 1773 2587 1787
rect 2613 1773 2627 1787
rect 2773 1773 2787 1787
rect 2813 1773 2827 1787
rect 2833 1773 2847 1787
rect 2873 1773 2887 1787
rect 3013 1773 3027 1787
rect 3053 1773 3067 1787
rect 3093 1773 3107 1787
rect 3173 1773 3187 1787
rect 3213 1773 3227 1787
rect 3313 1773 3327 1787
rect 3353 1773 3367 1787
rect 3513 1773 3527 1787
rect 3593 1773 3607 1787
rect 3633 1773 3647 1787
rect 3733 1773 3747 1787
rect 3773 1773 3787 1787
rect 3933 1773 3947 1787
rect 3973 1773 3987 1787
rect 4033 1773 4047 1787
rect 4073 1773 4087 1787
rect 4113 1773 4127 1787
rect 4313 1773 4327 1787
rect 4373 1773 4387 1787
rect 4413 1773 4427 1787
rect 4453 1773 4467 1787
rect 4533 1773 4547 1787
rect 4573 1773 4587 1787
rect 1073 1753 1087 1767
rect 1373 1753 1387 1767
rect 1613 1753 1627 1767
rect 2213 1753 2227 1767
rect 2253 1753 2267 1767
rect 2433 1753 2447 1767
rect 2513 1753 2527 1767
rect 2793 1753 2807 1767
rect 2933 1753 2947 1767
rect 3033 1753 3047 1767
rect 4093 1753 4107 1767
rect 4233 1753 4247 1767
rect 4273 1753 4287 1767
rect 4393 1753 4407 1767
rect 53 1613 67 1627
rect 133 1613 147 1627
rect 573 1613 587 1627
rect 713 1613 727 1627
rect 913 1613 927 1627
rect 1313 1613 1327 1627
rect 1433 1613 1447 1627
rect 1573 1613 1587 1627
rect 1913 1613 1927 1627
rect 1953 1613 1967 1627
rect 2213 1613 2227 1627
rect 2733 1613 2747 1627
rect 2813 1613 2827 1627
rect 2933 1613 2947 1627
rect 3013 1613 3027 1627
rect 3073 1613 3087 1627
rect 3693 1613 3707 1627
rect 3793 1613 3807 1627
rect 3933 1613 3947 1627
rect 4013 1613 4027 1627
rect 4073 1613 4087 1627
rect 4153 1613 4167 1627
rect 4253 1613 4267 1627
rect 4333 1613 4347 1627
rect 4413 1613 4427 1627
rect 4473 1613 4487 1627
rect 4573 1613 4587 1627
rect 93 1593 107 1607
rect 393 1593 407 1607
rect 433 1593 447 1607
rect 473 1593 487 1607
rect 513 1593 527 1607
rect 753 1593 767 1607
rect 953 1593 967 1607
rect 1133 1593 1147 1607
rect 1173 1593 1187 1607
rect 1353 1593 1367 1607
rect 1613 1593 1627 1607
rect 1753 1593 1767 1607
rect 1793 1593 1807 1607
rect 1873 1593 1887 1607
rect 2153 1593 2167 1607
rect 2193 1593 2207 1607
rect 2293 1593 2307 1607
rect 2373 1593 2387 1607
rect 2413 1593 2427 1607
rect 2553 1593 2567 1607
rect 2593 1593 2607 1607
rect 2633 1593 2647 1607
rect 2693 1593 2707 1607
rect 2713 1593 2727 1607
rect 2753 1593 2767 1607
rect 2853 1593 2867 1607
rect 2913 1593 2927 1607
rect 2953 1593 2967 1607
rect 3093 1593 3107 1607
rect 3133 1593 3147 1607
rect 3393 1593 3407 1607
rect 3433 1593 3447 1607
rect 3533 1593 3547 1607
rect 3573 1593 3587 1607
rect 3653 1593 3667 1607
rect 3853 1593 3867 1607
rect 3893 1593 3907 1607
rect 3913 1593 3927 1607
rect 3953 1593 3967 1607
rect 3993 1593 4007 1607
rect 4033 1593 4047 1607
rect 4193 1593 4207 1607
rect 4233 1593 4247 1607
rect 4273 1593 4287 1607
rect 4373 1593 4387 1607
rect 4593 1593 4607 1607
rect 4633 1593 4647 1607
rect 33 1573 47 1587
rect 113 1573 127 1587
rect 153 1573 167 1587
rect 173 1573 187 1587
rect 213 1573 227 1587
rect 293 1573 307 1587
rect 373 1573 387 1587
rect 413 1573 427 1587
rect 553 1573 567 1587
rect 593 1573 607 1587
rect 633 1573 647 1587
rect 693 1573 707 1587
rect 733 1573 747 1587
rect 793 1573 807 1587
rect 833 1573 847 1587
rect 893 1573 907 1587
rect 933 1573 947 1587
rect 993 1573 1007 1587
rect 1033 1573 1047 1587
rect 1113 1573 1127 1587
rect 1153 1573 1167 1587
rect 1193 1573 1207 1587
rect 1233 1573 1247 1587
rect 1293 1573 1307 1587
rect 1333 1573 1347 1587
rect 1413 1573 1427 1587
rect 1453 1573 1467 1587
rect 1493 1573 1507 1587
rect 1553 1573 1567 1587
rect 1593 1573 1607 1587
rect 1653 1573 1667 1587
rect 1693 1573 1707 1587
rect 1773 1573 1787 1587
rect 1813 1573 1827 1587
rect 1893 1573 1907 1587
rect 1933 1573 1947 1587
rect 1973 1573 1987 1587
rect 2013 1573 2027 1587
rect 2053 1573 2067 1587
rect 2133 1573 2147 1587
rect 2173 1573 2187 1587
rect 2233 1573 2247 1587
rect 2533 1573 2547 1587
rect 2573 1573 2587 1587
rect 2793 1573 2807 1587
rect 2833 1573 2847 1587
rect 2993 1573 3007 1587
rect 3053 1573 3067 1587
rect 3113 1573 3127 1587
rect 3153 1573 3167 1587
rect 3213 1573 3227 1587
rect 3313 1573 3327 1587
rect 3373 1573 3387 1587
rect 3413 1573 3427 1587
rect 3713 1573 3727 1587
rect 3773 1573 3787 1587
rect 3833 1573 3847 1587
rect 3873 1573 3887 1587
rect 4093 1573 4107 1587
rect 4133 1573 4147 1587
rect 4173 1573 4187 1587
rect 4313 1573 4327 1587
rect 4353 1573 4367 1587
rect 4433 1573 4447 1587
rect 4493 1573 4507 1587
rect 4553 1573 4567 1587
rect 4613 1573 4627 1587
rect 4653 1573 4667 1587
rect 4713 1573 4727 1587
rect 193 1553 207 1567
rect 233 1553 247 1567
rect 273 1553 287 1567
rect 313 1553 327 1567
rect 613 1553 627 1567
rect 653 1553 667 1567
rect 813 1553 827 1567
rect 853 1553 867 1567
rect 1013 1553 1027 1567
rect 1053 1553 1067 1567
rect 1213 1553 1227 1567
rect 1253 1553 1267 1567
rect 1473 1553 1487 1567
rect 1513 1553 1527 1567
rect 1673 1553 1687 1567
rect 1713 1553 1727 1567
rect 2033 1553 2047 1567
rect 2073 1553 2087 1567
rect 2653 1553 2667 1567
rect 3193 1553 3207 1567
rect 3233 1553 3247 1567
rect 3293 1553 3307 1567
rect 3333 1553 3347 1567
rect 4693 1553 4707 1567
rect 4733 1553 4747 1567
rect 133 1333 147 1347
rect 173 1333 187 1347
rect 233 1333 247 1347
rect 273 1333 287 1347
rect 333 1333 347 1347
rect 373 1333 387 1347
rect 833 1333 847 1347
rect 913 1333 927 1347
rect 953 1333 967 1347
rect 973 1333 987 1347
rect 1013 1333 1027 1347
rect 1073 1333 1087 1347
rect 1113 1333 1127 1347
rect 1253 1333 1267 1347
rect 1513 1333 1527 1347
rect 1553 1333 1567 1347
rect 1693 1333 1707 1347
rect 1733 1333 1747 1347
rect 1893 1333 1907 1347
rect 1933 1333 1947 1347
rect 2153 1333 2167 1347
rect 2193 1333 2207 1347
rect 2233 1333 2247 1347
rect 2273 1333 2287 1347
rect 2433 1333 2447 1347
rect 2473 1333 2487 1347
rect 4133 1333 4147 1347
rect 4173 1333 4187 1347
rect 4313 1333 4327 1347
rect 4353 1333 4367 1347
rect 53 1313 67 1327
rect 93 1313 107 1327
rect 113 1313 127 1327
rect 153 1313 167 1327
rect 213 1313 227 1327
rect 253 1313 267 1327
rect 353 1313 367 1327
rect 413 1313 427 1327
rect 453 1313 467 1327
rect 493 1313 507 1327
rect 533 1313 547 1327
rect 613 1313 627 1327
rect 653 1313 667 1327
rect 713 1313 727 1327
rect 753 1313 767 1327
rect 933 1313 947 1327
rect 993 1313 1007 1327
rect 1093 1313 1107 1327
rect 1133 1313 1147 1327
rect 1173 1313 1187 1327
rect 1333 1313 1347 1327
rect 1373 1313 1387 1327
rect 1433 1313 1447 1327
rect 1473 1313 1487 1327
rect 1533 1313 1547 1327
rect 1613 1313 1627 1327
rect 1653 1313 1667 1327
rect 1713 1313 1727 1327
rect 1773 1313 1787 1327
rect 1813 1313 1827 1327
rect 1873 1313 1887 1327
rect 1913 1313 1927 1327
rect 1993 1313 2007 1327
rect 2033 1313 2047 1327
rect 2093 1313 2107 1327
rect 2133 1313 2147 1327
rect 2173 1313 2187 1327
rect 2253 1313 2267 1327
rect 2373 1313 2387 1327
rect 2453 1313 2467 1327
rect 2513 1313 2527 1327
rect 2653 1313 2667 1327
rect 2693 1313 2707 1327
rect 2773 1313 2787 1327
rect 2813 1313 2827 1327
rect 3213 1313 3227 1327
rect 3253 1313 3267 1327
rect 3533 1313 3547 1327
rect 3753 1313 3767 1327
rect 4053 1313 4067 1327
rect 4093 1313 4107 1327
rect 4153 1313 4167 1327
rect 4333 1313 4347 1327
rect 4393 1313 4407 1327
rect 4433 1313 4447 1327
rect 4493 1313 4507 1327
rect 4533 1313 4547 1327
rect 4673 1313 4687 1327
rect 4733 1313 4747 1327
rect 33 1293 47 1307
rect 393 1293 407 1307
rect 433 1293 447 1307
rect 553 1293 567 1307
rect 593 1293 607 1307
rect 633 1293 647 1307
rect 693 1293 707 1307
rect 733 1293 747 1307
rect 793 1293 807 1307
rect 853 1293 867 1307
rect 1233 1293 1247 1307
rect 1293 1293 1307 1307
rect 1313 1293 1327 1307
rect 1353 1293 1367 1307
rect 1453 1293 1467 1307
rect 1493 1293 1507 1307
rect 1593 1293 1607 1307
rect 1633 1293 1647 1307
rect 1833 1293 1847 1307
rect 1973 1293 1987 1307
rect 2013 1293 2027 1307
rect 2333 1293 2347 1307
rect 2573 1293 2587 1307
rect 2613 1293 2627 1307
rect 2633 1293 2647 1307
rect 2673 1293 2687 1307
rect 2753 1293 2767 1307
rect 2793 1293 2807 1307
rect 2833 1293 2847 1307
rect 2933 1293 2947 1307
rect 2973 1293 2987 1307
rect 3053 1293 3067 1307
rect 3113 1293 3127 1307
rect 3153 1293 3167 1307
rect 3193 1293 3207 1307
rect 3353 1293 3367 1307
rect 3393 1293 3407 1307
rect 3473 1293 3487 1307
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3673 1293 3687 1307
rect 3713 1293 3727 1307
rect 3813 1293 3827 1307
rect 3893 1293 3907 1307
rect 3933 1293 3947 1307
rect 4033 1293 4047 1307
rect 4073 1293 4087 1307
rect 4233 1293 4247 1307
rect 4273 1293 4287 1307
rect 4413 1293 4427 1307
rect 4453 1293 4467 1307
rect 4513 1293 4527 1307
rect 4553 1293 4567 1307
rect 4573 1293 4587 1307
rect 4613 1293 4627 1307
rect 73 1273 87 1287
rect 513 1273 527 1287
rect 1193 1273 1207 1287
rect 1793 1273 1807 1287
rect 2073 1273 2087 1287
rect 2313 1273 2327 1287
rect 2493 1273 2507 1287
rect 3133 1273 3147 1287
rect 3233 1273 3247 1287
rect 3553 1273 3567 1287
rect 3613 1273 3627 1287
rect 3693 1273 3707 1287
rect 3733 1273 3747 1287
rect 4593 1273 4607 1287
rect 4653 1273 4667 1287
rect 4753 1273 4767 1287
rect 333 1133 347 1147
rect 533 1133 547 1147
rect 2353 1133 2367 1147
rect 2473 1133 2487 1147
rect 53 1113 67 1127
rect 93 1113 107 1127
rect 113 1113 127 1127
rect 153 1113 167 1127
rect 373 1113 387 1127
rect 573 1113 587 1127
rect 713 1113 727 1127
rect 773 1113 787 1127
rect 933 1113 947 1127
rect 973 1113 987 1127
rect 993 1113 1007 1127
rect 1033 1113 1047 1127
rect 1133 1113 1147 1127
rect 1173 1113 1187 1127
rect 1293 1113 1307 1127
rect 1353 1113 1367 1127
rect 1473 1113 1487 1127
rect 2053 1113 2067 1127
rect 2093 1113 2107 1127
rect 2133 1113 2147 1127
rect 2393 1113 2407 1127
rect 2593 1113 2607 1127
rect 2633 1113 2647 1127
rect 2673 1113 2687 1127
rect 2693 1113 2707 1127
rect 2733 1113 2747 1127
rect 2853 1113 2867 1127
rect 2893 1113 2907 1127
rect 2973 1113 2987 1127
rect 3133 1113 3147 1127
rect 3173 1113 3187 1127
rect 3213 1113 3227 1127
rect 3253 1113 3267 1127
rect 3333 1113 3347 1127
rect 3373 1113 3387 1127
rect 3393 1113 3407 1127
rect 3433 1113 3447 1127
rect 3873 1113 3887 1127
rect 3913 1113 3927 1127
rect 4053 1113 4067 1127
rect 4133 1113 4147 1127
rect 4173 1113 4187 1127
rect 4353 1113 4367 1127
rect 4393 1113 4407 1127
rect 4533 1113 4547 1127
rect 4573 1113 4587 1127
rect 33 1093 47 1107
rect 73 1093 87 1107
rect 133 1093 147 1107
rect 173 1093 187 1107
rect 213 1093 227 1107
rect 253 1093 267 1107
rect 313 1093 327 1107
rect 353 1093 367 1107
rect 413 1093 427 1107
rect 453 1093 467 1107
rect 513 1093 527 1107
rect 553 1093 567 1107
rect 653 1093 667 1107
rect 833 1093 847 1107
rect 873 1093 887 1107
rect 913 1093 927 1107
rect 953 1093 967 1107
rect 1013 1093 1027 1107
rect 1053 1093 1067 1107
rect 1113 1093 1127 1107
rect 1153 1093 1167 1107
rect 1233 1093 1247 1107
rect 1393 1093 1407 1107
rect 1493 1093 1507 1107
rect 1553 1093 1567 1107
rect 1633 1093 1647 1107
rect 1673 1093 1687 1107
rect 1713 1093 1727 1107
rect 1813 1093 1827 1107
rect 1853 1093 1867 1107
rect 1893 1093 1907 1107
rect 1973 1093 1987 1107
rect 2073 1093 2087 1107
rect 2113 1093 2127 1107
rect 2193 1093 2207 1107
rect 2233 1093 2247 1107
rect 2293 1093 2307 1107
rect 2333 1093 2347 1107
rect 2373 1093 2387 1107
rect 2453 1093 2467 1107
rect 2533 1093 2547 1107
rect 2613 1093 2627 1107
rect 2653 1093 2667 1107
rect 3033 1093 3047 1107
rect 3113 1093 3127 1107
rect 3153 1093 3167 1107
rect 3493 1093 3507 1107
rect 3633 1093 3647 1107
rect 3693 1093 3707 1107
rect 3833 1093 3847 1107
rect 3973 1093 3987 1107
rect 4293 1093 4307 1107
rect 4373 1093 4387 1107
rect 4413 1093 4427 1107
rect 4493 1093 4507 1107
rect 4553 1093 4567 1107
rect 4593 1093 4607 1107
rect 4633 1093 4647 1107
rect 4673 1093 4687 1107
rect 233 1073 247 1087
rect 273 1073 287 1087
rect 433 1073 447 1087
rect 473 1073 487 1087
rect 633 1073 647 1087
rect 673 1073 687 1087
rect 733 1073 747 1087
rect 813 1073 827 1087
rect 853 1073 867 1087
rect 1213 1073 1227 1087
rect 1253 1073 1267 1087
rect 1313 1073 1327 1087
rect 1373 1073 1387 1087
rect 1413 1073 1427 1087
rect 1533 1073 1547 1087
rect 1573 1073 1587 1087
rect 1613 1073 1627 1087
rect 1653 1073 1667 1087
rect 1693 1073 1707 1087
rect 1733 1073 1747 1087
rect 1793 1073 1807 1087
rect 1833 1073 1847 1087
rect 1873 1073 1887 1087
rect 1913 1073 1927 1087
rect 1953 1073 1967 1087
rect 1993 1073 2007 1087
rect 2173 1073 2187 1087
rect 2213 1073 2227 1087
rect 2273 1073 2287 1087
rect 2313 1073 2327 1087
rect 2513 1073 2527 1087
rect 2553 1073 2567 1087
rect 3013 1073 3027 1087
rect 3053 1073 3067 1087
rect 3953 1073 3967 1087
rect 3993 1073 4007 1087
rect 4273 1073 4287 1087
rect 4313 1073 4327 1087
rect 4473 1073 4487 1087
rect 4513 1073 4527 1087
rect 4653 1073 4667 1087
rect 4693 1073 4707 1087
rect 33 853 47 867
rect 73 853 87 867
rect 133 853 147 867
rect 733 853 747 867
rect 773 853 787 867
rect 853 853 867 867
rect 913 853 927 867
rect 953 853 967 867
rect 1013 853 1027 867
rect 1053 853 1067 867
rect 1213 853 1227 867
rect 1253 853 1267 867
rect 1473 853 1487 867
rect 1513 853 1527 867
rect 1533 853 1547 867
rect 1573 853 1587 867
rect 1753 853 1767 867
rect 1893 853 1907 867
rect 1933 853 1947 867
rect 2033 853 2047 867
rect 2073 853 2087 867
rect 2453 853 2467 867
rect 2493 853 2507 867
rect 2553 853 2567 867
rect 2593 853 2607 867
rect 2753 853 2767 867
rect 2793 853 2807 867
rect 3313 853 3327 867
rect 3353 853 3367 867
rect 53 833 67 847
rect 213 833 227 847
rect 253 833 267 847
rect 333 833 347 847
rect 373 833 387 847
rect 513 833 527 847
rect 573 833 587 847
rect 653 833 667 847
rect 693 833 707 847
rect 713 833 727 847
rect 753 833 767 847
rect 933 833 947 847
rect 1033 833 1047 847
rect 1073 833 1087 847
rect 1113 833 1127 847
rect 1153 833 1167 847
rect 1233 833 1247 847
rect 1273 833 1287 847
rect 1313 833 1327 847
rect 1373 833 1387 847
rect 1413 833 1427 847
rect 1493 833 1507 847
rect 1553 833 1567 847
rect 1633 833 1647 847
rect 1673 833 1687 847
rect 1833 833 1847 847
rect 1913 833 1927 847
rect 1973 833 1987 847
rect 2053 833 2067 847
rect 2093 833 2107 847
rect 2133 833 2147 847
rect 2193 833 2207 847
rect 2233 833 2247 847
rect 2313 833 2327 847
rect 2353 833 2367 847
rect 2393 833 2407 847
rect 2433 833 2447 847
rect 2473 833 2487 847
rect 2573 833 2587 847
rect 2613 833 2627 847
rect 2633 833 2647 847
rect 2673 833 2687 847
rect 2773 833 2787 847
rect 2853 833 2867 847
rect 2893 833 2907 847
rect 2953 833 2967 847
rect 3173 833 3187 847
rect 3233 833 3247 847
rect 3273 833 3287 847
rect 3333 833 3347 847
rect 3973 833 3987 847
rect 4013 833 4027 847
rect 4553 833 4567 847
rect 4593 833 4607 847
rect 4653 833 4667 847
rect 4693 833 4707 847
rect 113 813 127 827
rect 173 813 187 827
rect 233 813 247 827
rect 273 813 287 827
rect 313 813 327 827
rect 353 813 367 827
rect 393 813 407 827
rect 433 813 447 827
rect 473 813 487 827
rect 633 813 647 827
rect 833 813 847 827
rect 893 813 907 827
rect 1093 813 1107 827
rect 1133 813 1147 827
rect 1353 813 1367 827
rect 1393 813 1407 827
rect 1653 813 1667 827
rect 1693 813 1707 827
rect 1713 813 1727 827
rect 1773 813 1787 827
rect 2173 813 2187 827
rect 2213 813 2227 827
rect 2293 813 2307 827
rect 2693 813 2707 827
rect 2833 813 2847 827
rect 2873 813 2887 827
rect 2913 813 2927 827
rect 3013 813 3027 827
rect 3053 813 3067 827
rect 3093 813 3107 827
rect 3133 813 3147 827
rect 3213 813 3227 827
rect 3253 813 3267 827
rect 3413 813 3427 827
rect 3493 813 3507 827
rect 3533 813 3547 827
rect 3633 813 3647 827
rect 3673 813 3687 827
rect 3793 813 3807 827
rect 3833 813 3847 827
rect 3913 813 3927 827
rect 3993 813 4007 827
rect 4033 813 4047 827
rect 4073 813 4087 827
rect 4153 813 4167 827
rect 4193 813 4207 827
rect 4373 813 4387 827
rect 4413 813 4427 827
rect 4493 813 4507 827
rect 4533 813 4547 827
rect 4573 813 4587 827
rect 4633 813 4647 827
rect 4673 813 4687 827
rect 493 793 507 807
rect 593 793 607 807
rect 673 793 687 807
rect 1293 793 1307 807
rect 1853 793 1867 807
rect 1953 793 1967 807
rect 2113 793 2127 807
rect 2333 793 2347 807
rect 2373 793 2387 807
rect 2653 793 2667 807
rect 2973 793 2987 807
rect 3033 793 3047 807
rect 3113 793 3127 807
rect 3153 793 3167 807
rect 53 653 67 667
rect 153 653 167 667
rect 193 653 207 667
rect 313 653 327 667
rect 1193 653 1207 667
rect 1313 653 1327 667
rect 1593 653 1607 667
rect 1653 653 1667 667
rect 1993 653 2007 667
rect 2673 653 2687 667
rect 3133 653 3147 667
rect 3193 653 3207 667
rect 3393 653 3407 667
rect 33 633 47 647
rect 73 633 87 647
rect 113 633 127 647
rect 273 633 287 647
rect 493 633 507 647
rect 533 633 547 647
rect 573 633 587 647
rect 613 633 627 647
rect 673 633 687 647
rect 713 633 727 647
rect 753 633 767 647
rect 793 633 807 647
rect 813 633 827 647
rect 873 633 887 647
rect 913 633 927 647
rect 953 633 967 647
rect 1053 633 1067 647
rect 1093 633 1107 647
rect 1133 633 1147 647
rect 1233 633 1247 647
rect 1333 633 1347 647
rect 1373 633 1387 647
rect 1433 633 1447 647
rect 1473 633 1487 647
rect 1553 633 1567 647
rect 1693 633 1707 647
rect 1833 633 1847 647
rect 1873 633 1887 647
rect 1953 633 1967 647
rect 2033 633 2047 647
rect 2073 633 2087 647
rect 2273 633 2287 647
rect 2313 633 2327 647
rect 2333 633 2347 647
rect 2373 633 2387 647
rect 2873 633 2887 647
rect 2913 633 2927 647
rect 2993 633 3007 647
rect 3033 633 3047 647
rect 3073 633 3087 647
rect 3533 633 3547 647
rect 3573 633 3587 647
rect 3673 633 3687 647
rect 3713 633 3727 647
rect 3793 633 3807 647
rect 3833 633 3847 647
rect 3873 633 3887 647
rect 4033 633 4047 647
rect 4113 633 4127 647
rect 4153 633 4167 647
rect 4453 633 4467 647
rect 4493 633 4507 647
rect 4593 633 4607 647
rect 4633 633 4647 647
rect 4713 633 4727 647
rect 133 613 147 627
rect 173 613 187 627
rect 213 613 227 627
rect 293 613 307 627
rect 333 613 347 627
rect 353 613 367 627
rect 393 613 407 627
rect 473 613 487 627
rect 513 613 527 627
rect 653 613 667 627
rect 693 613 707 627
rect 933 613 947 627
rect 973 613 987 627
rect 1033 613 1047 627
rect 1073 613 1087 627
rect 1153 613 1167 627
rect 1173 613 1187 627
rect 1213 613 1227 627
rect 1293 613 1307 627
rect 1353 613 1367 627
rect 1393 613 1407 627
rect 1453 613 1467 627
rect 1493 613 1507 627
rect 1573 613 1587 627
rect 1613 613 1627 627
rect 1633 613 1647 627
rect 1673 613 1687 627
rect 1733 613 1747 627
rect 1773 613 1787 627
rect 1853 613 1867 627
rect 1893 613 1907 627
rect 1973 613 1987 627
rect 2013 613 2027 627
rect 2053 613 2067 627
rect 2093 613 2107 627
rect 2173 613 2187 627
rect 2213 613 2227 627
rect 2253 613 2267 627
rect 2293 613 2307 627
rect 2353 613 2367 627
rect 2393 613 2407 627
rect 2433 613 2447 627
rect 2473 613 2487 627
rect 2533 613 2547 627
rect 2573 613 2587 627
rect 2653 613 2667 627
rect 2693 613 2707 627
rect 2733 613 2747 627
rect 3053 613 3067 627
rect 3093 613 3107 627
rect 3153 613 3167 627
rect 3213 613 3227 627
rect 3253 613 3267 627
rect 3293 613 3307 627
rect 3373 613 3387 627
rect 3453 613 3467 627
rect 3513 613 3527 627
rect 3553 613 3567 627
rect 3853 613 3867 627
rect 3893 613 3907 627
rect 3973 613 3987 627
rect 4273 613 4287 627
rect 4353 613 4367 627
rect 4433 613 4447 627
rect 4473 613 4487 627
rect 373 593 387 607
rect 413 593 427 607
rect 853 593 867 607
rect 1753 593 1767 607
rect 1793 593 1807 607
rect 2153 593 2167 607
rect 2193 593 2207 607
rect 2453 593 2467 607
rect 2493 593 2507 607
rect 2553 593 2567 607
rect 2593 593 2607 607
rect 2713 593 2727 607
rect 2753 593 2767 607
rect 3273 593 3287 607
rect 3313 593 3327 607
rect 3433 593 3447 607
rect 3473 593 3487 607
rect 3953 593 3967 607
rect 3993 593 4007 607
rect 4253 593 4267 607
rect 4293 593 4307 607
rect 4333 593 4347 607
rect 4373 593 4387 607
rect 13 373 27 387
rect 53 373 67 387
rect 93 373 107 387
rect 133 373 147 387
rect 193 373 207 387
rect 233 373 247 387
rect 273 373 287 387
rect 313 373 327 387
rect 373 373 387 387
rect 453 373 467 387
rect 493 373 507 387
rect 533 373 547 387
rect 573 373 587 387
rect 833 373 847 387
rect 873 373 887 387
rect 893 373 907 387
rect 933 373 947 387
rect 993 373 1007 387
rect 1033 373 1047 387
rect 1073 373 1087 387
rect 1113 373 1127 387
rect 1773 373 1787 387
rect 1813 373 1827 387
rect 1953 373 1967 387
rect 1993 373 2007 387
rect 2033 373 2047 387
rect 2073 373 2087 387
rect 2113 373 2127 387
rect 2153 373 2167 387
rect 2293 373 2307 387
rect 2333 373 2347 387
rect 2453 373 2467 387
rect 2493 373 2507 387
rect 2613 373 2627 387
rect 2653 373 2667 387
rect 2893 373 2907 387
rect 2933 373 2947 387
rect 3673 373 3687 387
rect 3713 373 3727 387
rect 3753 373 3767 387
rect 3793 373 3807 387
rect 4313 373 4327 387
rect 4353 373 4367 387
rect 33 353 47 367
rect 113 353 127 367
rect 213 353 227 367
rect 293 353 307 367
rect 473 353 487 367
rect 553 353 567 367
rect 593 353 607 367
rect 653 353 667 367
rect 693 353 707 367
rect 853 353 867 367
rect 913 353 927 367
rect 1013 353 1027 367
rect 1093 353 1107 367
rect 1173 353 1187 367
rect 1213 353 1227 367
rect 1273 353 1287 367
rect 1313 353 1327 367
rect 1453 353 1467 367
rect 1493 353 1507 367
rect 1553 353 1567 367
rect 1633 353 1647 367
rect 1673 353 1687 367
rect 1713 353 1727 367
rect 1753 353 1767 367
rect 1793 353 1807 367
rect 1853 353 1867 367
rect 1893 353 1907 367
rect 1973 353 1987 367
rect 2053 353 2067 367
rect 2133 353 2147 367
rect 2313 353 2327 367
rect 2433 353 2447 367
rect 2473 353 2487 367
rect 2553 353 2567 367
rect 2633 353 2647 367
rect 2673 353 2687 367
rect 2693 353 2707 367
rect 2733 353 2747 367
rect 2913 353 2927 367
rect 2973 353 2987 367
rect 3013 353 3027 367
rect 3073 353 3087 367
rect 3113 353 3127 367
rect 3253 353 3267 367
rect 3313 353 3327 367
rect 3353 353 3367 367
rect 3433 353 3447 367
rect 3473 353 3487 367
rect 3633 353 3647 367
rect 3693 353 3707 367
rect 3773 353 3787 367
rect 3853 353 3867 367
rect 3893 353 3907 367
rect 3953 353 3967 367
rect 4013 353 4027 367
rect 4333 353 4347 367
rect 4393 353 4407 367
rect 4433 353 4447 367
rect 4493 353 4507 367
rect 353 333 367 347
rect 413 333 427 347
rect 633 333 647 347
rect 673 333 687 347
rect 713 333 727 347
rect 753 333 767 347
rect 793 333 807 347
rect 1153 333 1167 347
rect 1193 333 1207 347
rect 1233 333 1247 347
rect 1253 333 1267 347
rect 1293 333 1307 347
rect 1373 333 1387 347
rect 1413 333 1427 347
rect 1433 333 1447 347
rect 1473 333 1487 347
rect 1613 333 1627 347
rect 1913 333 1927 347
rect 2213 333 2227 347
rect 2253 333 2267 347
rect 2353 333 2367 347
rect 2393 333 2407 347
rect 2753 333 2767 347
rect 2793 333 2807 347
rect 2833 333 2847 347
rect 2993 333 3007 347
rect 3033 333 3047 347
rect 3093 333 3107 347
rect 3133 333 3147 347
rect 3173 333 3187 347
rect 3213 333 3227 347
rect 3333 333 3347 347
rect 3373 333 3387 347
rect 3413 333 3427 347
rect 3513 333 3527 347
rect 3553 333 3567 347
rect 3593 333 3607 347
rect 3873 333 3887 347
rect 3913 333 3927 347
rect 4073 333 4087 347
rect 4153 333 4167 347
rect 4193 333 4207 347
rect 4413 333 4427 347
rect 4453 333 4467 347
rect 4553 333 4567 347
rect 4633 333 4647 347
rect 4673 333 4687 347
rect 773 313 787 327
rect 1393 313 1407 327
rect 1533 313 1547 327
rect 1653 313 1667 327
rect 1693 313 1707 327
rect 1873 313 1887 327
rect 2233 313 2247 327
rect 2373 313 2387 327
rect 2573 313 2587 327
rect 2713 313 2727 327
rect 2813 313 2827 327
rect 3193 313 3207 327
rect 3273 313 3287 327
rect 3453 313 3467 327
rect 3533 313 3547 327
rect 3573 313 3587 327
rect 3973 313 3987 327
rect 4033 313 4047 327
rect 4513 313 4527 327
rect 133 173 147 187
rect 633 173 647 187
rect 773 173 787 187
rect 813 173 827 187
rect 1013 173 1027 187
rect 1493 173 1507 187
rect 1693 173 1707 187
rect 2553 173 2567 187
rect 2693 173 2707 187
rect 2853 173 2867 187
rect 3153 173 3167 187
rect 3253 173 3267 187
rect 3553 173 3567 187
rect 3833 173 3847 187
rect 4013 173 4027 187
rect 4093 173 4107 187
rect 4193 173 4207 187
rect 4453 173 4467 187
rect 4493 173 4507 187
rect 4673 173 4687 187
rect 173 153 187 167
rect 253 153 267 167
rect 293 153 307 167
rect 313 153 327 167
rect 353 153 367 167
rect 673 153 687 167
rect 733 153 747 167
rect 913 153 927 167
rect 953 153 967 167
rect 1033 153 1047 167
rect 1073 153 1087 167
rect 1133 153 1147 167
rect 1173 153 1187 167
rect 1453 153 1467 167
rect 1653 153 1667 167
rect 1913 153 1927 167
rect 1953 153 1967 167
rect 2013 153 2027 167
rect 2073 153 2087 167
rect 2093 153 2107 167
rect 2133 153 2147 167
rect 2273 153 2287 167
rect 2313 153 2327 167
rect 2353 153 2367 167
rect 2393 153 2407 167
rect 2433 153 2447 167
rect 2513 153 2527 167
rect 2593 153 2607 167
rect 2633 153 2647 167
rect 2993 153 3007 167
rect 3033 153 3047 167
rect 3113 153 3127 167
rect 3353 153 3367 167
rect 3393 153 3407 167
rect 3473 153 3487 167
rect 3533 153 3547 167
rect 3573 153 3587 167
rect 3613 153 3627 167
rect 3693 153 3707 167
rect 3733 153 3747 167
rect 3893 153 3907 167
rect 3933 153 3947 167
rect 3993 153 4007 167
rect 4033 153 4047 167
rect 4073 153 4087 167
rect 4113 153 4127 167
rect 4173 153 4187 167
rect 4213 153 4227 167
rect 4233 153 4247 167
rect 4273 153 4287 167
rect 4473 153 4487 167
rect 4513 153 4527 167
rect 53 133 67 147
rect 93 133 107 147
rect 113 133 127 147
rect 153 133 167 147
rect 233 133 247 147
rect 273 133 287 147
rect 333 133 347 147
rect 373 133 387 147
rect 453 133 467 147
rect 493 133 507 147
rect 513 133 527 147
rect 553 133 567 147
rect 613 133 627 147
rect 653 133 667 147
rect 753 133 767 147
rect 793 133 807 147
rect 833 133 847 147
rect 893 133 907 147
rect 933 133 947 147
rect 993 133 1007 147
rect 1053 133 1067 147
rect 1093 133 1107 147
rect 1153 133 1167 147
rect 1193 133 1207 147
rect 1233 133 1247 147
rect 1273 133 1287 147
rect 1333 133 1347 147
rect 1373 133 1387 147
rect 1473 133 1487 147
rect 1513 133 1527 147
rect 1533 133 1547 147
rect 1573 133 1587 147
rect 1673 133 1687 147
rect 1713 133 1727 147
rect 1733 133 1747 147
rect 1773 133 1787 147
rect 1853 133 1867 147
rect 2173 133 2187 147
rect 2213 133 2227 147
rect 2293 133 2307 147
rect 2333 133 2347 147
rect 2413 133 2427 147
rect 2453 133 2467 147
rect 2533 133 2547 147
rect 2573 133 2587 147
rect 2613 133 2627 147
rect 2653 133 2667 147
rect 2713 133 2727 147
rect 2753 133 2767 147
rect 2793 133 2807 147
rect 2873 133 2887 147
rect 3173 133 3187 147
rect 3233 133 3247 147
rect 3853 133 3867 147
rect 3913 133 3927 147
rect 3953 133 3967 147
rect 4253 133 4267 147
rect 4293 133 4307 147
rect 4373 133 4387 147
rect 4433 133 4447 147
rect 4573 133 4587 147
rect 4653 133 4667 147
rect 4713 133 4727 147
rect 33 113 47 127
rect 73 113 87 127
rect 433 113 447 127
rect 473 113 487 127
rect 533 113 547 127
rect 573 113 587 127
rect 1253 113 1267 127
rect 1293 113 1307 127
rect 1353 113 1367 127
rect 1393 113 1407 127
rect 1553 113 1567 127
rect 1593 113 1607 127
rect 1753 113 1767 127
rect 1793 113 1807 127
rect 1833 113 1847 127
rect 1873 113 1887 127
rect 2033 113 2047 127
rect 2193 113 2207 127
rect 2233 113 2247 127
rect 2773 113 2787 127
rect 2813 113 2827 127
rect 4353 113 4367 127
rect 4393 113 4407 127
rect 4553 113 4567 127
rect 4593 113 4607 127
rect 4693 113 4707 127
rect 4733 113 4747 127
<< labels >>
flabel metal1 s 4782 2 4842 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 1477 -23 1483 -17 7 FreeSans 16 270 0 0 Cin[5]
port 2 nsew
flabel metal2 s 1757 -23 1763 -17 7 FreeSans 16 270 0 0 Cin[4]
port 3 nsew
flabel metal2 s 1897 -23 1903 -17 7 FreeSans 16 270 0 0 Cin[3]
port 4 nsew
flabel metal2 s 1937 -23 1943 -17 7 FreeSans 16 270 0 0 Cin[2]
port 5 nsew
flabel metal2 s 1977 -23 1983 -17 7 FreeSans 16 270 0 0 Cin[1]
port 6 nsew
flabel metal2 s 2117 -23 2123 -17 7 FreeSans 16 270 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 3556 -16 3564 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal2 s 4077 4617 4083 4623 3 FreeSans 16 90 0 0 Vld
port 9 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 3476 -16 3484 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2756 -16 2764 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal2 s 4237 4617 4243 4623 3 FreeSans 16 90 0 0 Xout[3]
port 14 nsew
flabel metal2 s 4197 4617 4203 4623 3 FreeSans 16 90 0 0 Xout[2]
port 15 nsew
flabel metal2 s 4157 4617 4163 4623 3 FreeSans 16 90 0 0 Xout[1]
port 16 nsew
flabel metal2 s 4117 4617 4123 4623 3 FreeSans 16 90 0 0 Xout[0]
port 17 nsew
flabel metal3 s 4816 1316 4824 1324 3 FreeSans 16 0 0 0 Yin[3]
port 18 nsew
flabel metal3 s 4816 3676 4824 3684 3 FreeSans 16 0 0 0 Yin[2]
port 19 nsew
flabel metal3 s 4816 3716 4824 3724 3 FreeSans 16 0 0 0 Yin[1]
port 20 nsew
flabel metal3 s 4816 3956 4824 3964 3 FreeSans 16 0 0 0 Yin[0]
port 21 nsew
flabel metal2 s 4637 4617 4643 4623 3 FreeSans 16 90 0 0 Yout[3]
port 22 nsew
flabel metal2 s 4557 4617 4563 4623 3 FreeSans 16 90 0 0 Yout[2]
port 23 nsew
flabel metal2 s 4317 4617 4323 4623 3 FreeSans 16 90 0 0 Yout[1]
port 24 nsew
flabel metal2 s 4277 4617 4283 4623 3 FreeSans 16 90 0 0 Yout[0]
port 25 nsew
flabel metal2 s 4017 4617 4023 4623 3 FreeSans 16 90 0 0 clk
port 26 nsew
rlabel metal1 204 242 316 258 0 _989_.gnd
rlabel metal1 204 2 316 18 0 _989_.vdd
rlabel metal2 293 153 307 167 0 _989_.A
rlabel metal2 273 133 287 147 0 _989_.B
rlabel metal2 233 133 247 147 0 _989_.C
rlabel metal2 253 153 267 167 0 _989_.Y
rlabel metal1 164 242 256 258 0 _978_.gnd
rlabel metal1 164 482 256 498 0 _978_.vdd
rlabel metal2 233 373 247 387 0 _978_.A
rlabel metal2 193 373 207 387 0 _978_.B
rlabel metal2 213 353 227 367 0 _978_.Y
rlabel metal1 4 242 96 258 0 _975_.gnd
rlabel metal1 4 482 96 498 0 _975_.vdd
rlabel metal2 13 373 27 387 0 _975_.A
rlabel metal2 53 373 67 387 0 _975_.B
rlabel metal2 33 353 47 367 0 _975_.Y
rlabel metal1 84 242 176 258 0 _973_.gnd
rlabel metal1 84 482 176 498 0 _973_.vdd
rlabel metal2 93 373 107 387 0 _973_.A
rlabel metal2 133 373 147 387 0 _973_.B
rlabel metal2 113 353 127 367 0 _973_.Y
rlabel metal1 244 242 336 258 0 _971_.gnd
rlabel metal1 244 482 336 498 0 _971_.vdd
rlabel metal2 313 373 327 387 0 _971_.A
rlabel metal2 273 373 287 387 0 _971_.B
rlabel metal2 293 353 307 367 0 _971_.Y
rlabel metal1 104 242 216 258 0 _984_.gnd
rlabel metal1 104 2 216 18 0 _984_.vdd
rlabel metal2 113 133 127 147 0 _984_.A
rlabel metal2 133 173 147 187 0 _984_.B
rlabel metal2 153 133 167 147 0 _984_.C
rlabel metal2 173 153 187 167 0 _984_.Y
rlabel metal1 4 242 116 258 0 _976_.gnd
rlabel metal1 4 2 116 18 0 _976_.vdd
rlabel metal2 93 133 107 147 0 _976_.A
rlabel metal2 73 113 87 127 0 _976_.B
rlabel metal2 53 133 67 147 0 _976_.C
rlabel metal2 33 113 47 127 0 _976_.Y
rlabel metal1 304 242 416 258 0 _985_.gnd
rlabel metal1 304 2 416 18 0 _985_.vdd
rlabel metal2 313 153 327 167 0 _985_.A
rlabel metal2 333 133 347 147 0 _985_.B
rlabel metal2 373 133 387 147 0 _985_.C
rlabel metal2 353 153 367 167 0 _985_.Y
rlabel metal1 424 242 516 258 0 _925_.gnd
rlabel metal1 424 482 516 498 0 _925_.vdd
rlabel metal2 493 373 507 387 0 _925_.A
rlabel metal2 453 373 467 387 0 _925_.B
rlabel metal2 473 353 487 367 0 _925_.Y
rlabel metal1 404 242 516 258 0 _988_.gnd
rlabel metal1 404 2 516 18 0 _988_.vdd
rlabel metal2 493 133 507 147 0 _988_.A
rlabel metal2 473 113 487 127 0 _988_.B
rlabel metal2 453 133 467 147 0 _988_.C
rlabel metal2 433 113 447 127 0 _988_.Y
rlabel metal1 504 242 616 258 0 _986_.gnd
rlabel metal1 504 482 616 498 0 _986_.vdd
rlabel metal2 593 353 607 367 0 _986_.A
rlabel metal2 573 373 587 387 0 _986_.B
rlabel metal2 553 353 567 367 0 _986_.C
rlabel metal2 533 373 547 387 0 _986_.Y
rlabel metal1 504 242 616 258 0 _981_.gnd
rlabel metal1 504 2 616 18 0 _981_.vdd
rlabel metal2 513 133 527 147 0 _981_.A
rlabel metal2 533 113 547 127 0 _981_.B
rlabel metal2 553 133 567 147 0 _981_.C
rlabel metal2 573 113 587 127 0 _981_.Y
rlabel metal1 324 242 436 258 0 _918_.gnd
rlabel metal1 324 482 436 498 0 _918_.vdd
rlabel metal2 413 333 427 347 0 _918_.A
rlabel metal2 353 333 367 347 0 _918_.Y
rlabel metal2 373 373 387 387 0 _918_.B
rlabel metal1 604 242 716 258 0 _1050_.gnd
rlabel metal1 604 2 716 18 0 _1050_.vdd
rlabel metal2 613 133 627 147 0 _1050_.A
rlabel metal2 633 173 647 187 0 _1050_.B
rlabel metal2 653 133 667 147 0 _1050_.C
rlabel metal2 673 153 687 167 0 _1050_.Y
rlabel metal1 704 242 816 258 0 _970_.gnd
rlabel metal1 704 2 816 18 0 _970_.vdd
rlabel metal2 793 133 807 147 0 _970_.A
rlabel metal2 773 173 787 187 0 _970_.B
rlabel metal2 753 133 767 147 0 _970_.C
rlabel metal2 733 153 747 167 0 _970_.Y
rlabel metal1 724 242 816 258 0 _926_.gnd
rlabel metal1 724 482 816 498 0 _926_.vdd
rlabel metal2 753 333 767 347 0 _926_.B
rlabel metal2 793 333 807 347 0 _926_.A
rlabel metal2 773 313 787 327 0 _926_.Y
rlabel metal1 604 242 736 258 0 _920_.gnd
rlabel metal1 604 482 736 498 0 _920_.vdd
rlabel metal2 713 333 727 347 0 _920_.A
rlabel metal2 693 353 707 367 0 _920_.B
rlabel metal2 633 333 647 347 0 _920_.C
rlabel metal2 653 353 667 367 0 _920_.D
rlabel metal2 673 333 687 347 0 _920_.Y
rlabel metal1 864 242 976 258 0 _982_.gnd
rlabel metal1 864 2 976 18 0 _982_.vdd
rlabel metal2 953 153 967 167 0 _982_.A
rlabel metal2 933 133 947 147 0 _982_.B
rlabel metal2 893 133 907 147 0 _982_.C
rlabel metal2 913 153 927 167 0 _982_.Y
rlabel metal1 1024 242 1136 258 0 _927_.gnd
rlabel metal1 1024 2 1136 18 0 _927_.vdd
rlabel metal2 1033 153 1047 167 0 _927_.A
rlabel metal2 1053 133 1067 147 0 _927_.B
rlabel metal2 1093 133 1107 147 0 _927_.C
rlabel metal2 1073 153 1087 167 0 _927_.Y
rlabel metal1 1044 242 1136 258 0 _922_.gnd
rlabel metal1 1044 482 1136 498 0 _922_.vdd
rlabel metal2 1113 373 1127 387 0 _922_.A
rlabel metal2 1073 373 1087 387 0 _922_.B
rlabel metal2 1093 353 1107 367 0 _922_.Y
rlabel metal1 804 242 896 258 0 _919_.gnd
rlabel metal1 804 482 896 498 0 _919_.vdd
rlabel metal2 873 373 887 387 0 _919_.A
rlabel metal2 833 373 847 387 0 _919_.B
rlabel metal2 853 353 867 367 0 _919_.Y
rlabel metal1 964 242 1056 258 0 _891_.gnd
rlabel metal1 964 482 1056 498 0 _891_.vdd
rlabel metal2 1033 373 1047 387 0 _891_.A
rlabel metal2 993 373 1007 387 0 _891_.B
rlabel metal2 1013 353 1027 367 0 _891_.Y
rlabel metal1 884 242 976 258 0 _885_.gnd
rlabel metal1 884 482 976 498 0 _885_.vdd
rlabel metal2 893 373 907 387 0 _885_.A
rlabel metal2 933 373 947 387 0 _885_.B
rlabel metal2 913 353 927 367 0 _885_.Y
rlabel metal1 964 242 1036 258 0 _923_.gnd
rlabel metal1 964 2 1036 18 0 _923_.vdd
rlabel metal2 1013 173 1027 187 0 _923_.A
rlabel metal2 993 133 1007 147 0 _923_.Y
rlabel metal1 804 242 876 258 0 _921_.gnd
rlabel metal1 804 2 876 18 0 _921_.vdd
rlabel metal2 813 173 827 187 0 _921_.A
rlabel metal2 833 133 847 147 0 _921_.Y
rlabel metal1 1124 242 1236 258 0 _931_.gnd
rlabel metal1 1124 2 1236 18 0 _931_.vdd
rlabel metal2 1133 153 1147 167 0 _931_.A
rlabel metal2 1153 133 1167 147 0 _931_.B
rlabel metal2 1193 133 1207 147 0 _931_.C
rlabel metal2 1173 153 1187 167 0 _931_.Y
rlabel metal1 1244 242 1356 258 0 _917_.gnd
rlabel metal1 1244 482 1356 498 0 _917_.vdd
rlabel metal2 1253 333 1267 347 0 _917_.A
rlabel metal2 1273 353 1287 367 0 _917_.B
rlabel metal2 1313 353 1327 367 0 _917_.C
rlabel metal2 1293 333 1307 347 0 _917_.Y
rlabel metal1 1324 242 1436 258 0 _930_.gnd
rlabel metal1 1324 2 1436 18 0 _930_.vdd
rlabel metal2 1333 133 1347 147 0 _930_.A
rlabel metal2 1353 113 1367 127 0 _930_.B
rlabel metal2 1373 133 1387 147 0 _930_.C
rlabel metal2 1393 113 1407 127 0 _930_.Y
rlabel metal1 1224 242 1336 258 0 _924_.gnd
rlabel metal1 1224 2 1336 18 0 _924_.vdd
rlabel metal2 1233 133 1247 147 0 _924_.A
rlabel metal2 1253 113 1267 127 0 _924_.B
rlabel metal2 1273 133 1287 147 0 _924_.C
rlabel metal2 1293 113 1307 127 0 _924_.Y
rlabel metal1 1124 242 1256 258 0 _887_.gnd
rlabel metal1 1124 482 1256 498 0 _887_.vdd
rlabel metal2 1233 333 1247 347 0 _887_.A
rlabel metal2 1213 353 1227 367 0 _887_.B
rlabel metal2 1153 333 1167 347 0 _887_.C
rlabel metal2 1173 353 1187 367 0 _887_.D
rlabel metal2 1193 333 1207 347 0 _887_.Y
rlabel metal1 1424 242 1536 258 0 _888_.gnd
rlabel metal1 1424 482 1536 498 0 _888_.vdd
rlabel metal2 1433 333 1447 347 0 _888_.A
rlabel metal2 1453 353 1467 367 0 _888_.B
rlabel metal2 1493 353 1507 367 0 _888_.C
rlabel metal2 1473 333 1487 347 0 _888_.Y
rlabel metal1 1584 242 1696 258 0 _929_.gnd
rlabel metal1 1584 482 1696 498 0 _929_.vdd
rlabel metal2 1673 353 1687 367 0 _929_.A
rlabel metal2 1653 313 1667 327 0 _929_.B
rlabel metal2 1633 353 1647 367 0 _929_.C
rlabel metal2 1613 333 1627 347 0 _929_.Y
rlabel metal1 1424 242 1536 258 0 _928_.gnd
rlabel metal1 1424 2 1536 18 0 _928_.vdd
rlabel metal2 1513 133 1527 147 0 _928_.A
rlabel metal2 1493 173 1507 187 0 _928_.B
rlabel metal2 1473 133 1487 147 0 _928_.C
rlabel metal2 1453 153 1467 167 0 _928_.Y
rlabel metal1 1344 242 1436 258 0 _886_.gnd
rlabel metal1 1344 482 1436 498 0 _886_.vdd
rlabel metal2 1373 333 1387 347 0 _886_.B
rlabel metal2 1413 333 1427 347 0 _886_.A
rlabel metal2 1393 313 1407 327 0 _886_.Y
rlabel metal1 1524 242 1596 258 0 _892_.gnd
rlabel metal1 1524 482 1596 498 0 _892_.vdd
rlabel metal2 1533 313 1547 327 0 _892_.A
rlabel metal2 1553 353 1567 367 0 _892_.Y
rlabel metal1 1524 242 1636 258 0 _940_.gnd
rlabel metal1 1524 2 1636 18 0 _940_.vdd
rlabel metal2 1533 133 1547 147 0 _940_.A
rlabel metal2 1553 113 1567 127 0 _940_.B
rlabel metal2 1573 133 1587 147 0 _940_.C
rlabel metal2 1593 113 1607 127 0 _940_.Y
rlabel metal1 1824 242 1916 258 0 _884_.gnd
rlabel metal1 1824 2 1916 18 0 _884_.vdd
rlabel metal2 1833 113 1847 127 0 _884_.A
rlabel metal2 1873 113 1887 127 0 _884_.B
rlabel metal2 1853 133 1867 147 0 _884_.Y
rlabel metal1 1624 242 1736 258 0 _932_.gnd
rlabel metal1 1624 2 1736 18 0 _932_.vdd
rlabel metal2 1713 133 1727 147 0 _932_.A
rlabel metal2 1693 173 1707 187 0 _932_.B
rlabel metal2 1673 133 1687 147 0 _932_.C
rlabel metal2 1653 153 1667 167 0 _932_.Y
rlabel metal1 1844 242 1956 258 0 _896_.gnd
rlabel metal1 1844 482 1956 498 0 _896_.vdd
rlabel metal2 1853 353 1867 367 0 _896_.A
rlabel metal2 1873 313 1887 327 0 _896_.B
rlabel metal2 1893 353 1907 367 0 _896_.C
rlabel metal2 1913 333 1927 347 0 _896_.Y
rlabel metal1 1684 242 1756 258 0 _889_.gnd
rlabel metal1 1684 482 1756 498 0 _889_.vdd
rlabel metal2 1693 313 1707 327 0 _889_.A
rlabel metal2 1713 353 1727 367 0 _889_.Y
rlabel metal1 1724 242 1836 258 0 _939_.gnd
rlabel metal1 1724 2 1836 18 0 _939_.vdd
rlabel metal2 1733 133 1747 147 0 _939_.A
rlabel metal2 1753 113 1767 127 0 _939_.B
rlabel metal2 1773 133 1787 147 0 _939_.C
rlabel metal2 1793 113 1807 127 0 _939_.Y
rlabel metal1 1744 242 1856 258 0 _893_.gnd
rlabel metal1 1744 482 1856 498 0 _893_.vdd
rlabel metal2 1753 353 1767 367 0 _893_.A
rlabel metal2 1773 373 1787 387 0 _893_.B
rlabel metal2 1793 353 1807 367 0 _893_.C
rlabel metal2 1813 373 1827 387 0 _893_.Y
rlabel metal1 1904 242 1996 258 0 BUFX2_insert30.gnd
rlabel metal1 1904 2 1996 18 0 BUFX2_insert30.vdd
rlabel metal2 1913 153 1927 167 0 BUFX2_insert30.A
rlabel metal2 1953 153 1967 167 0 BUFX2_insert30.Y
rlabel metal1 2084 242 2176 258 0 BUFX2_insert23.gnd
rlabel metal1 2084 2 2176 18 0 BUFX2_insert23.vdd
rlabel metal2 2093 153 2107 167 0 BUFX2_insert23.A
rlabel metal2 2133 153 2147 167 0 BUFX2_insert23.Y
rlabel metal1 2024 242 2116 258 0 _866_.gnd
rlabel metal1 2024 482 2116 498 0 _866_.vdd
rlabel metal2 2033 373 2047 387 0 _866_.A
rlabel metal2 2073 373 2087 387 0 _866_.B
rlabel metal2 2053 353 2067 367 0 _866_.Y
rlabel metal1 1944 242 2036 258 0 _865_.gnd
rlabel metal1 1944 482 2036 498 0 _865_.vdd
rlabel metal2 1953 373 1967 387 0 _865_.A
rlabel metal2 1993 373 2007 387 0 _865_.B
rlabel metal2 1973 353 1987 367 0 _865_.Y
rlabel metal1 2104 242 2196 258 0 _856_.gnd
rlabel metal1 2104 482 2196 498 0 _856_.vdd
rlabel metal2 2113 373 2127 387 0 _856_.A
rlabel metal2 2153 373 2167 387 0 _856_.B
rlabel metal2 2133 353 2147 367 0 _856_.Y
rlabel metal1 1984 242 2096 258 0 _871_.gnd
rlabel metal1 1984 2 2096 18 0 _871_.vdd
rlabel metal2 2073 153 2087 167 0 _871_.A
rlabel metal2 2013 153 2027 167 0 _871_.Y
rlabel metal2 2033 113 2047 127 0 _871_.B
rlabel metal1 2384 242 2496 258 0 _895_.gnd
rlabel metal1 2384 2 2496 18 0 _895_.vdd
rlabel metal2 2393 153 2407 167 0 _895_.A
rlabel metal2 2413 133 2427 147 0 _895_.B
rlabel metal2 2453 133 2467 147 0 _895_.C
rlabel metal2 2433 153 2447 167 0 _895_.Y
rlabel metal1 2264 242 2356 258 0 _855_.gnd
rlabel metal1 2264 482 2356 498 0 _855_.vdd
rlabel metal2 2333 373 2347 387 0 _855_.A
rlabel metal2 2293 373 2307 387 0 _855_.B
rlabel metal2 2313 353 2327 367 0 _855_.Y
rlabel metal1 2184 242 2276 258 0 _867_.gnd
rlabel metal1 2184 482 2276 498 0 _867_.vdd
rlabel metal2 2213 333 2227 347 0 _867_.B
rlabel metal2 2253 333 2267 347 0 _867_.A
rlabel metal2 2233 313 2247 327 0 _867_.Y
rlabel metal1 2344 242 2436 258 0 _857_.gnd
rlabel metal1 2344 482 2436 498 0 _857_.vdd
rlabel metal2 2393 333 2407 347 0 _857_.B
rlabel metal2 2353 333 2367 347 0 _857_.A
rlabel metal2 2373 313 2387 327 0 _857_.Y
rlabel metal1 2164 242 2276 258 0 _872_.gnd
rlabel metal1 2164 2 2276 18 0 _872_.vdd
rlabel metal2 2173 133 2187 147 0 _872_.A
rlabel metal2 2193 113 2207 127 0 _872_.B
rlabel metal2 2213 133 2227 147 0 _872_.C
rlabel metal2 2233 113 2247 127 0 _872_.Y
rlabel metal1 2264 242 2396 258 0 _868_.gnd
rlabel metal1 2264 2 2396 18 0 _868_.vdd
rlabel metal2 2273 153 2287 167 0 _868_.A
rlabel metal2 2293 133 2307 147 0 _868_.B
rlabel metal2 2353 153 2367 167 0 _868_.C
rlabel metal2 2333 133 2347 147 0 _868_.D
rlabel metal2 2313 153 2327 167 0 _868_.Y
rlabel metal1 2584 242 2696 258 0 _869_.gnd
rlabel metal1 2584 2 2696 18 0 _869_.vdd
rlabel metal2 2593 153 2607 167 0 _869_.A
rlabel metal2 2613 133 2627 147 0 _869_.B
rlabel metal2 2653 133 2667 147 0 _869_.C
rlabel metal2 2633 153 2647 167 0 _869_.Y
rlabel metal1 2484 242 2596 258 0 _883_.gnd
rlabel metal1 2484 2 2596 18 0 _883_.vdd
rlabel metal2 2573 133 2587 147 0 _883_.A
rlabel metal2 2553 173 2567 187 0 _883_.B
rlabel metal2 2533 133 2547 147 0 _883_.C
rlabel metal2 2513 153 2527 167 0 _883_.Y
rlabel metal1 2524 242 2596 258 0 _876_.gnd
rlabel metal1 2524 482 2596 498 0 _876_.vdd
rlabel metal2 2573 313 2587 327 0 _876_.A
rlabel metal2 2553 353 2567 367 0 _876_.Y
rlabel metal1 2584 242 2696 258 0 _875_.gnd
rlabel metal1 2584 482 2696 498 0 _875_.vdd
rlabel metal2 2673 353 2687 367 0 _875_.A
rlabel metal2 2653 373 2667 387 0 _875_.B
rlabel metal2 2633 353 2647 367 0 _875_.C
rlabel metal2 2613 373 2627 387 0 _875_.Y
rlabel metal1 2424 242 2536 258 0 _852_.gnd
rlabel metal1 2424 482 2536 498 0 _852_.vdd
rlabel metal2 2433 353 2447 367 0 _852_.A
rlabel metal2 2453 373 2467 387 0 _852_.B
rlabel metal2 2473 353 2487 367 0 _852_.C
rlabel metal2 2493 373 2507 387 0 _852_.Y
rlabel metal1 2904 242 3156 258 0 _1546_.gnd
rlabel metal1 2904 2 3156 18 0 _1546_.vdd
rlabel metal2 2993 153 3007 167 0 _1546_.D
rlabel metal2 3033 153 3047 167 0 _1546_.CLK
rlabel metal2 3113 153 3127 167 0 _1546_.Q
rlabel metal1 2864 242 2956 258 0 _879_.gnd
rlabel metal1 2864 482 2956 498 0 _879_.vdd
rlabel metal2 2933 373 2947 387 0 _879_.A
rlabel metal2 2893 373 2907 387 0 _879_.B
rlabel metal2 2913 353 2927 367 0 _879_.Y
rlabel metal1 2684 242 2796 258 0 _877_.gnd
rlabel metal1 2684 482 2796 498 0 _877_.vdd
rlabel metal2 2693 353 2707 367 0 _877_.A
rlabel metal2 2713 313 2727 327 0 _877_.B
rlabel metal2 2733 353 2747 367 0 _877_.C
rlabel metal2 2753 333 2767 347 0 _877_.Y
rlabel metal1 2784 242 2876 258 0 _878_.gnd
rlabel metal1 2784 482 2876 498 0 _878_.vdd
rlabel metal2 2833 333 2847 347 0 _878_.B
rlabel metal2 2793 333 2807 347 0 _878_.A
rlabel metal2 2813 313 2827 327 0 _878_.Y
rlabel metal1 2844 242 2916 258 0 _873_.gnd
rlabel metal1 2844 2 2916 18 0 _873_.vdd
rlabel metal2 2853 173 2867 187 0 _873_.A
rlabel metal2 2873 133 2887 147 0 _873_.Y
rlabel metal1 2684 242 2756 258 0 _870_.gnd
rlabel metal1 2684 2 2756 18 0 _870_.vdd
rlabel metal2 2693 173 2707 187 0 _870_.A
rlabel metal2 2713 133 2727 147 0 _870_.Y
rlabel metal1 2744 242 2856 258 0 _874_.gnd
rlabel metal1 2744 2 2856 18 0 _874_.vdd
rlabel metal2 2753 133 2767 147 0 _874_.A
rlabel metal2 2773 113 2787 127 0 _874_.B
rlabel metal2 2793 133 2807 147 0 _874_.C
rlabel metal2 2813 113 2827 127 0 _874_.Y
rlabel metal1 3044 242 3156 258 0 _880_.gnd
rlabel metal1 3044 482 3156 498 0 _880_.vdd
rlabel metal2 3133 333 3147 347 0 _880_.A
rlabel metal2 3113 353 3127 367 0 _880_.B
rlabel metal2 3073 353 3087 367 0 _880_.C
rlabel metal2 3093 333 3107 347 0 _880_.Y
rlabel metal1 2944 242 3056 258 0 _853_.gnd
rlabel metal1 2944 482 3056 498 0 _853_.vdd
rlabel metal2 3033 333 3047 347 0 _853_.A
rlabel metal2 3013 353 3027 367 0 _853_.B
rlabel metal2 2973 353 2987 367 0 _853_.C
rlabel metal2 2993 333 3007 347 0 _853_.Y
rlabel metal1 3144 242 3236 258 0 _1334_.gnd
rlabel metal1 3144 482 3236 498 0 _1334_.vdd
rlabel metal2 3173 333 3187 347 0 _1334_.B
rlabel metal2 3213 333 3227 347 0 _1334_.A
rlabel metal2 3193 313 3207 327 0 _1334_.Y
rlabel metal1 3204 242 3276 258 0 _864_.gnd
rlabel metal1 3204 2 3276 18 0 _864_.vdd
rlabel metal2 3253 173 3267 187 0 _864_.A
rlabel metal2 3233 133 3247 147 0 _864_.Y
rlabel metal1 3144 242 3216 258 0 _851_.gnd
rlabel metal1 3144 2 3216 18 0 _851_.vdd
rlabel metal2 3153 173 3167 187 0 _851_.A
rlabel metal2 3173 133 3187 147 0 _851_.Y
rlabel metal1 3264 242 3516 258 0 _1548_.gnd
rlabel metal1 3264 2 3516 18 0 _1548_.vdd
rlabel metal2 3353 153 3367 167 0 _1548_.D
rlabel metal2 3393 153 3407 167 0 _1548_.CLK
rlabel metal2 3473 153 3487 167 0 _1548_.Q
rlabel metal1 3284 242 3396 258 0 _811_.gnd
rlabel metal1 3284 482 3396 498 0 _811_.vdd
rlabel metal2 3373 333 3387 347 0 _811_.A
rlabel metal2 3353 353 3367 367 0 _811_.B
rlabel metal2 3313 353 3327 367 0 _811_.C
rlabel metal2 3333 333 3347 347 0 _811_.Y
rlabel metal1 3384 242 3496 258 0 _1341_.gnd
rlabel metal1 3384 482 3496 498 0 _1341_.vdd
rlabel metal2 3473 353 3487 367 0 _1341_.A
rlabel metal2 3453 313 3467 327 0 _1341_.B
rlabel metal2 3433 353 3447 367 0 _1341_.C
rlabel metal2 3413 333 3427 347 0 _1341_.Y
rlabel metal1 3224 242 3296 258 0 _809_.gnd
rlabel metal1 3224 482 3296 498 0 _809_.vdd
rlabel metal2 3273 313 3287 327 0 _809_.A
rlabel metal2 3253 353 3267 367 0 _809_.Y
rlabel metal1 3584 242 3836 258 0 _1532_.gnd
rlabel metal1 3584 2 3836 18 0 _1532_.vdd
rlabel metal2 3733 153 3747 167 0 _1532_.D
rlabel metal2 3693 153 3707 167 0 _1532_.CLK
rlabel metal2 3613 153 3627 167 0 _1532_.Q
rlabel metal1 3664 242 3756 258 0 _1336_.gnd
rlabel metal1 3664 482 3756 498 0 _1336_.vdd
rlabel metal2 3673 373 3687 387 0 _1336_.A
rlabel metal2 3713 373 3727 387 0 _1336_.B
rlabel metal2 3693 353 3707 367 0 _1336_.Y
rlabel metal1 3484 242 3576 258 0 _1335_.gnd
rlabel metal1 3484 482 3576 498 0 _1335_.vdd
rlabel metal2 3513 333 3527 347 0 _1335_.B
rlabel metal2 3553 333 3567 347 0 _1335_.A
rlabel metal2 3533 313 3547 327 0 _1335_.Y
rlabel metal1 3504 242 3596 258 0 _1333_.gnd
rlabel metal1 3504 2 3596 18 0 _1333_.vdd
rlabel metal2 3533 153 3547 167 0 _1333_.B
rlabel metal2 3573 153 3587 167 0 _1333_.A
rlabel metal2 3553 173 3567 187 0 _1333_.Y
rlabel metal1 3564 242 3676 258 0 _1337_.gnd
rlabel metal1 3564 482 3676 498 0 _1337_.vdd
rlabel metal2 3573 313 3587 327 0 _1337_.A
rlabel metal2 3593 333 3607 347 0 _1337_.B
rlabel metal2 3633 353 3647 367 0 _1337_.Y
rlabel metal1 3884 242 3996 258 0 _1332_.gnd
rlabel metal1 3884 2 3996 18 0 _1332_.vdd
rlabel metal2 3893 153 3907 167 0 _1332_.A
rlabel metal2 3913 133 3927 147 0 _1332_.B
rlabel metal2 3953 133 3967 147 0 _1332_.C
rlabel metal2 3933 153 3947 167 0 _1332_.Y
rlabel metal1 3824 242 3936 258 0 _863_.gnd
rlabel metal1 3824 482 3936 498 0 _863_.vdd
rlabel metal2 3913 333 3927 347 0 _863_.A
rlabel metal2 3893 353 3907 367 0 _863_.B
rlabel metal2 3853 353 3867 367 0 _863_.C
rlabel metal2 3873 333 3887 347 0 _863_.Y
rlabel metal1 3744 242 3836 258 0 _1338_.gnd
rlabel metal1 3744 482 3836 498 0 _1338_.vdd
rlabel metal2 3753 373 3767 387 0 _1338_.A
rlabel metal2 3793 373 3807 387 0 _1338_.B
rlabel metal2 3773 353 3787 367 0 _1338_.Y
rlabel metal1 3984 242 4076 258 0 _1324_.gnd
rlabel metal1 3984 2 4076 18 0 _1324_.vdd
rlabel metal2 4033 153 4047 167 0 _1324_.B
rlabel metal2 3993 153 4007 167 0 _1324_.A
rlabel metal2 4013 173 4027 187 0 _1324_.Y
rlabel metal1 3924 242 3996 258 0 _854_.gnd
rlabel metal1 3924 482 3996 498 0 _854_.vdd
rlabel metal2 3973 313 3987 327 0 _854_.A
rlabel metal2 3953 353 3967 367 0 _854_.Y
rlabel metal1 3824 242 3896 258 0 _806_.gnd
rlabel metal1 3824 2 3896 18 0 _806_.vdd
rlabel metal2 3833 173 3847 187 0 _806_.A
rlabel metal2 3853 133 3867 147 0 _806_.Y
rlabel metal1 3984 242 4056 258 0 _778_.gnd
rlabel metal1 3984 482 4056 498 0 _778_.vdd
rlabel metal2 4033 313 4047 327 0 _778_.A
rlabel metal2 4013 353 4027 367 0 _778_.Y
rlabel metal1 4044 242 4296 258 0 _1547_.gnd
rlabel metal1 4044 482 4296 498 0 _1547_.vdd
rlabel metal2 4193 333 4207 347 0 _1547_.D
rlabel metal2 4153 333 4167 347 0 _1547_.CLK
rlabel metal2 4073 333 4087 347 0 _1547_.Q
rlabel metal1 4224 242 4336 258 0 _1328_.gnd
rlabel metal1 4224 2 4336 18 0 _1328_.vdd
rlabel metal2 4233 153 4247 167 0 _1328_.A
rlabel metal2 4253 133 4267 147 0 _1328_.B
rlabel metal2 4293 133 4307 147 0 _1328_.C
rlabel metal2 4273 153 4287 167 0 _1328_.Y
rlabel metal1 4144 242 4236 258 0 _1326_.gnd
rlabel metal1 4144 2 4236 18 0 _1326_.vdd
rlabel metal2 4173 153 4187 167 0 _1326_.B
rlabel metal2 4213 153 4227 167 0 _1326_.A
rlabel metal2 4193 173 4207 187 0 _1326_.Y
rlabel metal1 4064 242 4156 258 0 _1325_.gnd
rlabel metal1 4064 2 4156 18 0 _1325_.vdd
rlabel metal2 4113 153 4127 167 0 _1325_.B
rlabel metal2 4073 153 4087 167 0 _1325_.A
rlabel metal2 4093 173 4107 187 0 _1325_.Y
rlabel metal1 4524 242 4776 258 0 _1530_.gnd
rlabel metal1 4524 482 4776 498 0 _1530_.vdd
rlabel metal2 4673 333 4687 347 0 _1530_.D
rlabel metal2 4633 333 4647 347 0 _1530_.CLK
rlabel metal2 4553 333 4567 347 0 _1530_.Q
rlabel metal1 4364 242 4476 258 0 _805_.gnd
rlabel metal1 4364 482 4476 498 0 _805_.vdd
rlabel metal2 4453 333 4467 347 0 _805_.A
rlabel metal2 4433 353 4447 367 0 _805_.B
rlabel metal2 4393 353 4407 367 0 _805_.C
rlabel metal2 4413 333 4427 347 0 _805_.Y
rlabel metal1 4284 242 4376 258 0 _1329_.gnd
rlabel metal1 4284 482 4376 498 0 _1329_.vdd
rlabel metal2 4353 373 4367 387 0 _1329_.A
rlabel metal2 4313 373 4327 387 0 _1329_.B
rlabel metal2 4333 353 4347 367 0 _1329_.Y
rlabel metal1 4324 242 4416 258 0 _1327_.gnd
rlabel metal1 4324 2 4416 18 0 _1327_.vdd
rlabel metal2 4393 113 4407 127 0 _1327_.A
rlabel metal2 4353 113 4367 127 0 _1327_.B
rlabel metal2 4373 133 4387 147 0 _1327_.Y
rlabel metal1 4464 242 4556 258 0 _1318_.gnd
rlabel metal1 4464 2 4556 18 0 _1318_.vdd
rlabel metal2 4513 153 4527 167 0 _1318_.B
rlabel metal2 4473 153 4487 167 0 _1318_.A
rlabel metal2 4493 173 4507 187 0 _1318_.Y
rlabel metal1 4404 242 4476 258 0 _1319_.gnd
rlabel metal1 4404 2 4476 18 0 _1319_.vdd
rlabel metal2 4453 173 4467 187 0 _1319_.A
rlabel metal2 4433 133 4447 147 0 _1319_.Y
rlabel metal1 4464 242 4536 258 0 _803_.gnd
rlabel metal1 4464 482 4536 498 0 _803_.vdd
rlabel metal2 4513 313 4527 327 0 _803_.A
rlabel metal2 4493 353 4507 367 0 _803_.Y
rlabel metal1 4684 242 4776 258 0 _1321_.gnd
rlabel metal1 4684 2 4776 18 0 _1321_.vdd
rlabel metal2 4693 113 4707 127 0 _1321_.A
rlabel metal2 4733 113 4747 127 0 _1321_.B
rlabel metal2 4713 133 4727 147 0 _1321_.Y
rlabel metal1 4544 242 4636 258 0 _1320_.gnd
rlabel metal1 4544 2 4636 18 0 _1320_.vdd
rlabel metal2 4553 113 4567 127 0 _1320_.A
rlabel metal2 4593 113 4607 127 0 _1320_.B
rlabel metal2 4573 133 4587 147 0 _1320_.Y
rlabel metal1 4624 242 4696 258 0 _848_.gnd
rlabel metal1 4624 2 4696 18 0 _848_.vdd
rlabel metal2 4673 173 4687 187 0 _848_.A
rlabel metal2 4653 133 4667 147 0 _848_.Y
rlabel metal1 84 722 196 738 0 _1026_.gnd
rlabel metal1 84 482 196 498 0 _1026_.vdd
rlabel metal2 173 613 187 627 0 _1026_.A
rlabel metal2 153 653 167 667 0 _1026_.B
rlabel metal2 133 613 147 627 0 _1026_.C
rlabel metal2 113 633 127 647 0 _1026_.Y
rlabel metal1 244 722 356 738 0 _983_.gnd
rlabel metal1 244 482 356 498 0 _983_.vdd
rlabel metal2 333 613 347 627 0 _983_.A
rlabel metal2 313 653 327 667 0 _983_.B
rlabel metal2 293 613 307 627 0 _983_.C
rlabel metal2 273 633 287 647 0 _983_.Y
rlabel metal1 4 722 96 738 0 _1025_.gnd
rlabel metal1 4 482 96 498 0 _1025_.vdd
rlabel metal2 33 633 47 647 0 _1025_.B
rlabel metal2 73 633 87 647 0 _1025_.A
rlabel metal2 53 653 67 667 0 _1025_.Y
rlabel metal1 184 722 256 738 0 _977_.gnd
rlabel metal1 184 482 256 498 0 _977_.vdd
rlabel metal2 193 653 207 667 0 _977_.A
rlabel metal2 213 613 227 627 0 _977_.Y
rlabel metal1 444 722 556 738 0 _979_.gnd
rlabel metal1 444 482 556 498 0 _979_.vdd
rlabel metal2 533 633 547 647 0 _979_.A
rlabel metal2 513 613 527 627 0 _979_.B
rlabel metal2 473 613 487 627 0 _979_.C
rlabel metal2 493 633 507 647 0 _979_.Y
rlabel metal1 344 722 456 738 0 _980_.gnd
rlabel metal1 344 482 456 498 0 _980_.vdd
rlabel metal2 353 613 367 627 0 _980_.A
rlabel metal2 373 593 387 607 0 _980_.B
rlabel metal2 393 613 407 627 0 _980_.C
rlabel metal2 413 593 427 607 0 _980_.Y
rlabel metal1 544 722 636 738 0 BUFX2_insert32.gnd
rlabel metal1 544 482 636 498 0 BUFX2_insert32.vdd
rlabel metal2 613 633 627 647 0 BUFX2_insert32.A
rlabel metal2 573 633 587 647 0 BUFX2_insert32.Y
rlabel metal1 724 722 816 738 0 BUFX2_insert24.gnd
rlabel metal1 724 482 816 498 0 BUFX2_insert24.vdd
rlabel metal2 793 633 807 647 0 BUFX2_insert24.A
rlabel metal2 753 633 767 647 0 BUFX2_insert24.Y
rlabel metal1 624 722 736 738 0 _1051_.gnd
rlabel metal1 624 482 736 498 0 _1051_.vdd
rlabel metal2 713 633 727 647 0 _1051_.A
rlabel metal2 693 613 707 627 0 _1051_.B
rlabel metal2 653 613 667 627 0 _1051_.C
rlabel metal2 673 633 687 647 0 _1051_.Y
rlabel metal1 904 722 1016 738 0 _901_.gnd
rlabel metal1 904 482 1016 498 0 _901_.vdd
rlabel metal2 913 633 927 647 0 _901_.A
rlabel metal2 933 613 947 627 0 _901_.B
rlabel metal2 973 613 987 627 0 _901_.C
rlabel metal2 953 633 967 647 0 _901_.Y
rlabel metal1 1004 722 1116 738 0 _898_.gnd
rlabel metal1 1004 482 1116 498 0 _898_.vdd
rlabel metal2 1093 633 1107 647 0 _898_.A
rlabel metal2 1073 613 1087 627 0 _898_.B
rlabel metal2 1033 613 1047 627 0 _898_.C
rlabel metal2 1053 633 1067 647 0 _898_.Y
rlabel metal1 804 722 916 738 0 _890_.gnd
rlabel metal1 804 482 916 498 0 _890_.vdd
rlabel metal2 813 633 827 647 0 _890_.A
rlabel metal2 873 633 887 647 0 _890_.Y
rlabel metal2 853 593 867 607 0 _890_.B
rlabel metal1 1324 722 1436 738 0 _992_.gnd
rlabel metal1 1324 482 1436 498 0 _992_.vdd
rlabel metal2 1333 633 1347 647 0 _992_.A
rlabel metal2 1353 613 1367 627 0 _992_.B
rlabel metal2 1393 613 1407 627 0 _992_.C
rlabel metal2 1373 633 1387 647 0 _992_.Y
rlabel metal1 1164 722 1276 738 0 _902_.gnd
rlabel metal1 1164 482 1276 498 0 _902_.vdd
rlabel metal2 1173 613 1187 627 0 _902_.A
rlabel metal2 1193 653 1207 667 0 _902_.B
rlabel metal2 1213 613 1227 627 0 _902_.C
rlabel metal2 1233 633 1247 647 0 _902_.Y
rlabel metal1 1264 722 1336 738 0 _941_.gnd
rlabel metal1 1264 482 1336 498 0 _941_.vdd
rlabel metal2 1313 653 1327 667 0 _941_.A
rlabel metal2 1293 613 1307 627 0 _941_.Y
rlabel metal1 1104 722 1176 738 0 _897_.gnd
rlabel metal1 1104 482 1176 498 0 _897_.vdd
rlabel metal2 1153 613 1167 627 0 _897_.A
rlabel metal2 1133 633 1147 647 0 _897_.Y
rlabel metal1 1424 722 1536 738 0 _938_.gnd
rlabel metal1 1424 482 1536 498 0 _938_.vdd
rlabel metal2 1433 633 1447 647 0 _938_.A
rlabel metal2 1453 613 1467 627 0 _938_.B
rlabel metal2 1493 613 1507 627 0 _938_.C
rlabel metal2 1473 633 1487 647 0 _938_.Y
rlabel metal1 1524 722 1636 738 0 _957_.gnd
rlabel metal1 1524 482 1636 498 0 _957_.vdd
rlabel metal2 1613 613 1627 627 0 _957_.A
rlabel metal2 1593 653 1607 667 0 _957_.B
rlabel metal2 1573 613 1587 627 0 _957_.C
rlabel metal2 1553 633 1567 647 0 _957_.Y
rlabel metal1 1824 722 1936 738 0 _861_.gnd
rlabel metal1 1824 482 1936 498 0 _861_.vdd
rlabel metal2 1833 633 1847 647 0 _861_.A
rlabel metal2 1853 613 1867 627 0 _861_.B
rlabel metal2 1893 613 1907 627 0 _861_.C
rlabel metal2 1873 633 1887 647 0 _861_.Y
rlabel metal1 1624 722 1736 738 0 _946_.gnd
rlabel metal1 1624 482 1736 498 0 _946_.vdd
rlabel metal2 1633 613 1647 627 0 _946_.A
rlabel metal2 1653 653 1667 667 0 _946_.B
rlabel metal2 1673 613 1687 627 0 _946_.C
rlabel metal2 1693 633 1707 647 0 _946_.Y
rlabel metal1 1724 722 1836 738 0 _942_.gnd
rlabel metal1 1724 482 1836 498 0 _942_.vdd
rlabel metal2 1733 613 1747 627 0 _942_.A
rlabel metal2 1753 593 1767 607 0 _942_.B
rlabel metal2 1773 613 1787 627 0 _942_.C
rlabel metal2 1793 593 1807 607 0 _942_.Y
rlabel metal1 2024 722 2136 738 0 _916_.gnd
rlabel metal1 2024 482 2136 498 0 _916_.vdd
rlabel metal2 2033 633 2047 647 0 _916_.A
rlabel metal2 2053 613 2067 627 0 _916_.B
rlabel metal2 2093 613 2107 627 0 _916_.C
rlabel metal2 2073 633 2087 647 0 _916_.Y
rlabel metal1 1924 722 2036 738 0 _915_.gnd
rlabel metal1 1924 482 2036 498 0 _915_.vdd
rlabel metal2 2013 613 2027 627 0 _915_.A
rlabel metal2 1993 653 2007 667 0 _915_.B
rlabel metal2 1973 613 1987 627 0 _915_.C
rlabel metal2 1953 633 1967 647 0 _915_.Y
rlabel metal1 2124 722 2236 738 0 _906_.gnd
rlabel metal1 2124 482 2236 498 0 _906_.vdd
rlabel metal2 2213 613 2227 627 0 _906_.A
rlabel metal2 2193 593 2207 607 0 _906_.B
rlabel metal2 2173 613 2187 627 0 _906_.C
rlabel metal2 2153 593 2167 607 0 _906_.Y
rlabel metal1 2324 722 2436 738 0 _907_.gnd
rlabel metal1 2324 482 2436 498 0 _907_.vdd
rlabel metal2 2333 633 2347 647 0 _907_.A
rlabel metal2 2353 613 2367 627 0 _907_.B
rlabel metal2 2393 613 2407 627 0 _907_.C
rlabel metal2 2373 633 2387 647 0 _907_.Y
rlabel metal1 2224 722 2336 738 0 _903_.gnd
rlabel metal1 2224 482 2336 498 0 _903_.vdd
rlabel metal2 2313 633 2327 647 0 _903_.A
rlabel metal2 2293 613 2307 627 0 _903_.B
rlabel metal2 2253 613 2267 627 0 _903_.C
rlabel metal2 2273 633 2287 647 0 _903_.Y
rlabel metal1 2624 722 2696 738 0 _858_.gnd
rlabel metal1 2624 482 2696 498 0 _858_.vdd
rlabel metal2 2673 653 2687 667 0 _858_.A
rlabel metal2 2653 613 2667 627 0 _858_.Y
rlabel metal1 2524 722 2636 738 0 _904_.gnd
rlabel metal1 2524 482 2636 498 0 _904_.vdd
rlabel metal2 2533 613 2547 627 0 _904_.A
rlabel metal2 2553 593 2567 607 0 _904_.B
rlabel metal2 2573 613 2587 627 0 _904_.C
rlabel metal2 2593 593 2607 607 0 _904_.Y
rlabel metal1 2424 722 2536 738 0 _894_.gnd
rlabel metal1 2424 482 2536 498 0 _894_.vdd
rlabel metal2 2433 613 2447 627 0 _894_.A
rlabel metal2 2453 593 2467 607 0 _894_.B
rlabel metal2 2473 613 2487 627 0 _894_.C
rlabel metal2 2493 593 2507 607 0 _894_.Y
rlabel metal1 2784 722 3036 738 0 _1549_.gnd
rlabel metal1 2784 482 3036 498 0 _1549_.vdd
rlabel metal2 2873 633 2887 647 0 _1549_.D
rlabel metal2 2913 633 2927 647 0 _1549_.CLK
rlabel metal2 2993 633 3007 647 0 _1549_.Q
rlabel metal1 2684 722 2796 738 0 _862_.gnd
rlabel metal1 2684 482 2796 498 0 _862_.vdd
rlabel metal2 2693 613 2707 627 0 _862_.A
rlabel metal2 2713 593 2727 607 0 _862_.B
rlabel metal2 2733 613 2747 627 0 _862_.C
rlabel metal2 2753 593 2767 607 0 _862_.Y
rlabel metal1 3024 722 3136 738 0 _1355_.gnd
rlabel metal1 3024 482 3136 498 0 _1355_.vdd
rlabel metal2 3033 633 3047 647 0 _1355_.A
rlabel metal2 3053 613 3067 627 0 _1355_.B
rlabel metal2 3093 613 3107 627 0 _1355_.C
rlabel metal2 3073 633 3087 647 0 _1355_.Y
rlabel metal1 3124 722 3196 738 0 _1347_.gnd
rlabel metal1 3124 482 3196 498 0 _1347_.vdd
rlabel metal2 3133 653 3147 667 0 _1347_.A
rlabel metal2 3153 613 3167 627 0 _1347_.Y
rlabel metal1 3184 722 3256 738 0 _1346_.gnd
rlabel metal1 3184 482 3256 498 0 _1346_.vdd
rlabel metal2 3193 653 3207 667 0 _1346_.A
rlabel metal2 3213 613 3227 627 0 _1346_.Y
rlabel metal1 3404 722 3496 738 0 _807_.gnd
rlabel metal1 3404 482 3496 498 0 _807_.vdd
rlabel metal2 3473 593 3487 607 0 _807_.A
rlabel metal2 3433 593 3447 607 0 _807_.B
rlabel metal2 3453 613 3467 627 0 _807_.Y
rlabel metal1 3344 722 3416 738 0 _1345_.gnd
rlabel metal1 3344 482 3416 498 0 _1345_.vdd
rlabel metal2 3393 653 3407 667 0 _1345_.A
rlabel metal2 3373 613 3387 627 0 _1345_.Y
rlabel metal1 3244 722 3356 738 0 _1348_.gnd
rlabel metal1 3244 482 3356 498 0 _1348_.vdd
rlabel metal2 3253 613 3267 627 0 _1348_.A
rlabel metal2 3273 593 3287 607 0 _1348_.B
rlabel metal2 3293 613 3307 627 0 _1348_.C
rlabel metal2 3313 593 3327 607 0 _1348_.Y
rlabel metal1 3584 722 3836 738 0 _1531_.gnd
rlabel metal1 3584 482 3836 498 0 _1531_.vdd
rlabel metal2 3673 633 3687 647 0 _1531_.D
rlabel metal2 3713 633 3727 647 0 _1531_.CLK
rlabel metal2 3793 633 3807 647 0 _1531_.Q
rlabel metal1 3484 722 3596 738 0 _808_.gnd
rlabel metal1 3484 482 3596 498 0 _808_.vdd
rlabel metal2 3573 633 3587 647 0 _808_.A
rlabel metal2 3553 613 3567 627 0 _808_.B
rlabel metal2 3513 613 3527 627 0 _808_.C
rlabel metal2 3533 633 3547 647 0 _808_.Y
rlabel metal1 4004 722 4256 738 0 _1562_.gnd
rlabel metal1 4004 482 4256 498 0 _1562_.vdd
rlabel metal2 4153 633 4167 647 0 _1562_.D
rlabel metal2 4113 633 4127 647 0 _1562_.CLK
rlabel metal2 4033 633 4047 647 0 _1562_.Q
rlabel metal1 3824 722 3936 738 0 _1340_.gnd
rlabel metal1 3824 482 3936 498 0 _1340_.vdd
rlabel metal2 3833 633 3847 647 0 _1340_.A
rlabel metal2 3853 613 3867 627 0 _1340_.B
rlabel metal2 3893 613 3907 627 0 _1340_.C
rlabel metal2 3873 633 3887 647 0 _1340_.Y
rlabel metal1 3924 722 4016 738 0 _1339_.gnd
rlabel metal1 3924 482 4016 498 0 _1339_.vdd
rlabel metal2 3993 593 4007 607 0 _1339_.A
rlabel metal2 3953 593 3967 607 0 _1339_.B
rlabel metal2 3973 613 3987 627 0 _1339_.Y
rlabel metal1 4244 722 4336 738 0 _804_.gnd
rlabel metal1 4244 482 4336 498 0 _804_.vdd
rlabel metal2 4253 593 4267 607 0 _804_.A
rlabel metal2 4293 593 4307 607 0 _804_.B
rlabel metal2 4273 613 4287 627 0 _804_.Y
rlabel metal1 4504 722 4756 738 0 _1545_.gnd
rlabel metal1 4504 482 4756 498 0 _1545_.vdd
rlabel metal2 4593 633 4607 647 0 _1545_.D
rlabel metal2 4633 633 4647 647 0 _1545_.CLK
rlabel metal2 4713 633 4727 647 0 _1545_.Q
rlabel metal1 4404 722 4516 738 0 _1323_.gnd
rlabel metal1 4404 482 4516 498 0 _1323_.vdd
rlabel metal2 4493 633 4507 647 0 _1323_.A
rlabel metal2 4473 613 4487 627 0 _1323_.B
rlabel metal2 4433 613 4447 627 0 _1323_.C
rlabel metal2 4453 633 4467 647 0 _1323_.Y
rlabel metal1 4324 722 4416 738 0 _1322_.gnd
rlabel metal1 4324 482 4416 498 0 _1322_.vdd
rlabel metal2 4333 593 4347 607 0 _1322_.A
rlabel metal2 4373 593 4387 607 0 _1322_.B
rlabel metal2 4353 613 4367 627 0 _1322_.Y
rlabel nsubstratencontact 4764 492 4764 492 0 FILL71250x7350.vdd
rlabel metal1 4744 722 4776 738 0 FILL71250x7350.gnd
rlabel metal1 184 722 296 738 0 _1040_.gnd
rlabel metal1 184 962 296 978 0 _1040_.vdd
rlabel metal2 273 813 287 827 0 _1040_.A
rlabel metal2 253 833 267 847 0 _1040_.B
rlabel metal2 213 833 227 847 0 _1040_.C
rlabel metal2 233 813 247 827 0 _1040_.Y
rlabel metal1 4 722 96 738 0 _974_.gnd
rlabel metal1 4 962 96 978 0 _974_.vdd
rlabel metal2 73 853 87 867 0 _974_.A
rlabel metal2 33 853 47 867 0 _974_.B
rlabel metal2 53 833 67 847 0 _974_.Y
rlabel metal1 84 722 196 738 0 _972_.gnd
rlabel metal1 84 962 196 978 0 _972_.vdd
rlabel metal2 173 813 187 827 0 _972_.A
rlabel metal2 113 813 127 827 0 _972_.Y
rlabel metal2 133 853 147 867 0 _972_.B
rlabel metal1 404 722 496 738 0 BUFX2_insert22.gnd
rlabel metal1 404 962 496 978 0 BUFX2_insert22.vdd
rlabel metal2 473 813 487 827 0 BUFX2_insert22.A
rlabel metal2 433 813 447 827 0 BUFX2_insert22.Y
rlabel metal1 484 722 556 738 0 _900_.gnd
rlabel metal1 484 962 556 978 0 _900_.vdd
rlabel metal2 493 793 507 807 0 _900_.A
rlabel metal2 513 833 527 847 0 _900_.Y
rlabel metal1 284 722 416 738 0 _1039_.gnd
rlabel metal1 284 962 416 978 0 _1039_.vdd
rlabel metal2 393 813 407 827 0 _1039_.A
rlabel metal2 373 833 387 847 0 _1039_.B
rlabel metal2 313 813 327 827 0 _1039_.C
rlabel metal2 333 833 347 847 0 _1039_.D
rlabel metal2 353 813 367 827 0 _1039_.Y
rlabel metal1 604 722 716 738 0 _1013_.gnd
rlabel metal1 604 962 716 978 0 _1013_.vdd
rlabel metal2 693 833 707 847 0 _1013_.A
rlabel metal2 673 793 687 807 0 _1013_.B
rlabel metal2 653 833 667 847 0 _1013_.C
rlabel metal2 633 813 647 827 0 _1013_.Y
rlabel metal1 544 722 616 738 0 _1012_.gnd
rlabel metal1 544 962 616 978 0 _1012_.vdd
rlabel metal2 593 793 607 807 0 _1012_.A
rlabel metal2 573 833 587 847 0 _1012_.Y
rlabel metal1 704 722 816 738 0 _990_.gnd
rlabel metal1 704 962 816 978 0 _990_.vdd
rlabel metal2 713 833 727 847 0 _990_.A
rlabel metal2 733 853 747 867 0 _990_.B
rlabel metal2 753 833 767 847 0 _990_.C
rlabel metal2 773 853 787 867 0 _990_.Y
rlabel metal1 904 722 996 738 0 _969_.gnd
rlabel metal1 904 962 996 978 0 _969_.vdd
rlabel metal2 913 853 927 867 0 _969_.A
rlabel metal2 953 853 967 867 0 _969_.B
rlabel metal2 933 833 947 847 0 _969_.Y
rlabel metal1 984 722 1096 738 0 _964_.gnd
rlabel metal1 984 962 1096 978 0 _964_.vdd
rlabel metal2 1073 833 1087 847 0 _964_.A
rlabel metal2 1053 853 1067 867 0 _964_.B
rlabel metal2 1033 833 1047 847 0 _964_.C
rlabel metal2 1013 853 1027 867 0 _964_.Y
rlabel metal1 804 722 916 738 0 _987_.gnd
rlabel metal1 804 962 916 978 0 _987_.vdd
rlabel metal2 893 813 907 827 0 _987_.A
rlabel metal2 833 813 847 827 0 _987_.Y
rlabel metal2 853 853 867 867 0 _987_.B
rlabel metal1 1084 722 1196 738 0 _963_.gnd
rlabel metal1 1084 962 1196 978 0 _963_.vdd
rlabel metal2 1093 813 1107 827 0 _963_.A
rlabel metal2 1113 833 1127 847 0 _963_.B
rlabel metal2 1153 833 1167 847 0 _963_.C
rlabel metal2 1133 813 1147 827 0 _963_.Y
rlabel metal1 1284 722 1356 738 0 _965_.gnd
rlabel metal1 1284 962 1356 978 0 _965_.vdd
rlabel metal2 1293 793 1307 807 0 _965_.A
rlabel metal2 1313 833 1327 847 0 _965_.Y
rlabel metal1 1184 722 1296 738 0 _968_.gnd
rlabel metal1 1184 962 1296 978 0 _968_.vdd
rlabel metal2 1273 833 1287 847 0 _968_.A
rlabel metal2 1253 853 1267 867 0 _968_.B
rlabel metal2 1233 833 1247 847 0 _968_.C
rlabel metal2 1213 853 1227 867 0 _968_.Y
rlabel metal1 1344 722 1456 738 0 _967_.gnd
rlabel metal1 1344 962 1456 978 0 _967_.vdd
rlabel metal2 1353 813 1367 827 0 _967_.A
rlabel metal2 1373 833 1387 847 0 _967_.B
rlabel metal2 1413 833 1427 847 0 _967_.C
rlabel metal2 1393 813 1407 827 0 _967_.Y
rlabel metal1 1604 722 1716 738 0 _937_.gnd
rlabel metal1 1604 962 1716 978 0 _937_.vdd
rlabel metal2 1693 813 1707 827 0 _937_.A
rlabel metal2 1673 833 1687 847 0 _937_.B
rlabel metal2 1633 833 1647 847 0 _937_.C
rlabel metal2 1653 813 1667 827 0 _937_.Y
rlabel metal1 1444 722 1536 738 0 _958_.gnd
rlabel metal1 1444 962 1536 978 0 _958_.vdd
rlabel metal2 1513 853 1527 867 0 _958_.A
rlabel metal2 1473 853 1487 867 0 _958_.B
rlabel metal2 1493 833 1507 847 0 _958_.Y
rlabel metal1 1524 722 1616 738 0 _933_.gnd
rlabel metal1 1524 962 1616 978 0 _933_.vdd
rlabel metal2 1533 853 1547 867 0 _933_.A
rlabel metal2 1573 853 1587 867 0 _933_.B
rlabel metal2 1553 833 1567 847 0 _933_.Y
rlabel metal1 1864 722 1956 738 0 _882_.gnd
rlabel metal1 1864 962 1956 978 0 _882_.vdd
rlabel metal2 1933 853 1947 867 0 _882_.A
rlabel metal2 1893 853 1907 867 0 _882_.B
rlabel metal2 1913 833 1927 847 0 _882_.Y
rlabel metal1 1804 722 1876 738 0 _859_.gnd
rlabel metal1 1804 962 1876 978 0 _859_.vdd
rlabel metal2 1853 793 1867 807 0 _859_.A
rlabel metal2 1833 833 1847 847 0 _859_.Y
rlabel metal1 1704 722 1816 738 0 _954_.gnd
rlabel metal1 1704 962 1816 978 0 _954_.vdd
rlabel metal2 1713 813 1727 827 0 _954_.A
rlabel metal2 1773 813 1787 827 0 _954_.Y
rlabel metal2 1753 853 1767 867 0 _954_.B
rlabel metal1 2104 722 2176 738 0 _947_.gnd
rlabel metal1 2104 962 2176 978 0 _947_.vdd
rlabel metal2 2113 793 2127 807 0 _947_.A
rlabel metal2 2133 833 2147 847 0 _947_.Y
rlabel metal1 1944 722 2016 738 0 _905_.gnd
rlabel metal1 1944 962 2016 978 0 _905_.vdd
rlabel metal2 1953 793 1967 807 0 _905_.A
rlabel metal2 1973 833 1987 847 0 _905_.Y
rlabel metal1 2004 722 2116 738 0 _943_.gnd
rlabel metal1 2004 962 2116 978 0 _943_.vdd
rlabel metal2 2093 833 2107 847 0 _943_.A
rlabel metal2 2073 853 2087 867 0 _943_.B
rlabel metal2 2053 833 2067 847 0 _943_.C
rlabel metal2 2033 853 2047 867 0 _943_.Y
rlabel metal1 2164 722 2276 738 0 _948_.gnd
rlabel metal1 2164 962 2276 978 0 _948_.vdd
rlabel metal2 2173 813 2187 827 0 _948_.A
rlabel metal2 2193 833 2207 847 0 _948_.B
rlabel metal2 2233 833 2247 847 0 _948_.C
rlabel metal2 2213 813 2227 827 0 _948_.Y
rlabel metal1 2264 722 2376 738 0 _945_.gnd
rlabel metal1 2264 962 2376 978 0 _945_.vdd
rlabel metal2 2353 833 2367 847 0 _945_.A
rlabel metal2 2333 793 2347 807 0 _945_.B
rlabel metal2 2313 833 2327 847 0 _945_.C
rlabel metal2 2293 813 2307 827 0 _945_.Y
rlabel metal1 2364 722 2436 738 0 _944_.gnd
rlabel metal1 2364 962 2436 978 0 _944_.vdd
rlabel metal2 2373 793 2387 807 0 _944_.A
rlabel metal2 2393 833 2407 847 0 _944_.Y
rlabel metal1 2624 722 2736 738 0 _909_.gnd
rlabel metal1 2624 962 2736 978 0 _909_.vdd
rlabel metal2 2633 833 2647 847 0 _909_.A
rlabel metal2 2653 793 2667 807 0 _909_.B
rlabel metal2 2673 833 2687 847 0 _909_.C
rlabel metal2 2693 813 2707 827 0 _909_.Y
rlabel metal1 2524 722 2636 738 0 _910_.gnd
rlabel metal1 2524 962 2636 978 0 _910_.vdd
rlabel metal2 2613 833 2627 847 0 _910_.A
rlabel metal2 2593 853 2607 867 0 _910_.B
rlabel metal2 2573 833 2587 847 0 _910_.C
rlabel metal2 2553 853 2567 867 0 _910_.Y
rlabel metal1 2424 722 2536 738 0 _908_.gnd
rlabel metal1 2424 962 2536 978 0 _908_.vdd
rlabel metal2 2433 833 2447 847 0 _908_.A
rlabel metal2 2453 853 2467 867 0 _908_.B
rlabel metal2 2473 833 2487 847 0 _908_.C
rlabel metal2 2493 853 2507 867 0 _908_.Y
rlabel metal1 2724 722 2816 738 0 _911_.gnd
rlabel metal1 2724 962 2816 978 0 _911_.vdd
rlabel metal2 2793 853 2807 867 0 _911_.A
rlabel metal2 2753 853 2767 867 0 _911_.B
rlabel metal2 2773 833 2787 847 0 _911_.Y
rlabel metal1 2924 722 2996 738 0 _881_.gnd
rlabel metal1 2924 962 2996 978 0 _881_.vdd
rlabel metal2 2973 793 2987 807 0 _881_.A
rlabel metal2 2953 833 2967 847 0 _881_.Y
rlabel metal1 2804 722 2936 738 0 _912_.gnd
rlabel metal1 2804 962 2936 978 0 _912_.vdd
rlabel metal2 2913 813 2927 827 0 _912_.A
rlabel metal2 2893 833 2907 847 0 _912_.B
rlabel metal2 2833 813 2847 827 0 _912_.C
rlabel metal2 2873 813 2887 827 0 _912_.Y
rlabel metal2 2853 833 2867 847 0 _912_.D
rlabel metal1 3204 722 3316 738 0 _1344_.gnd
rlabel metal1 3204 962 3316 978 0 _1344_.vdd
rlabel metal2 3213 813 3227 827 0 _1344_.A
rlabel metal2 3233 833 3247 847 0 _1344_.B
rlabel metal2 3273 833 3287 847 0 _1344_.C
rlabel metal2 3253 813 3267 827 0 _1344_.Y
rlabel metal1 3064 722 3156 738 0 _1343_.gnd
rlabel metal1 3064 962 3156 978 0 _1343_.vdd
rlabel metal2 3093 813 3107 827 0 _1343_.B
rlabel metal2 3133 813 3147 827 0 _1343_.A
rlabel metal2 3113 793 3127 807 0 _1343_.Y
rlabel metal1 2984 722 3076 738 0 _1342_.gnd
rlabel metal1 2984 962 3076 978 0 _1342_.vdd
rlabel metal2 3013 813 3027 827 0 _1342_.B
rlabel metal2 3053 813 3067 827 0 _1342_.A
rlabel metal2 3033 793 3047 807 0 _1342_.Y
rlabel metal1 3144 722 3216 738 0 _812_.gnd
rlabel metal1 3144 962 3216 978 0 _812_.vdd
rlabel metal2 3153 793 3167 807 0 _812_.A
rlabel metal2 3173 833 3187 847 0 _812_.Y
rlabel metal1 3384 722 3636 738 0 _1533_.gnd
rlabel metal1 3384 962 3636 978 0 _1533_.vdd
rlabel metal2 3533 813 3547 827 0 _1533_.D
rlabel metal2 3493 813 3507 827 0 _1533_.CLK
rlabel metal2 3413 813 3427 827 0 _1533_.Q
rlabel metal1 3304 722 3396 738 0 _1349_.gnd
rlabel metal1 3304 962 3396 978 0 _1349_.vdd
rlabel metal2 3313 853 3327 867 0 _1349_.A
rlabel metal2 3353 853 3367 867 0 _1349_.B
rlabel metal2 3333 833 3347 847 0 _1349_.Y
rlabel metal1 3624 722 3716 738 0 BUFX2_insert18.gnd
rlabel metal1 3624 962 3716 978 0 BUFX2_insert18.vdd
rlabel metal2 3633 813 3647 827 0 BUFX2_insert18.A
rlabel metal2 3673 813 3687 827 0 BUFX2_insert18.Y
rlabel metal1 3704 722 3956 738 0 _1561_.gnd
rlabel metal1 3704 962 3956 978 0 _1561_.vdd
rlabel metal2 3793 813 3807 827 0 _1561_.D
rlabel metal2 3833 813 3847 827 0 _1561_.CLK
rlabel metal2 3913 813 3927 827 0 _1561_.Q
rlabel metal1 3944 722 4056 738 0 _1331_.gnd
rlabel metal1 3944 962 4056 978 0 _1331_.vdd
rlabel metal2 4033 813 4047 827 0 _1331_.A
rlabel metal2 4013 833 4027 847 0 _1331_.B
rlabel metal2 3973 833 3987 847 0 _1331_.C
rlabel metal2 3993 813 4007 827 0 _1331_.Y
rlabel metal1 4044 722 4296 738 0 _1560_.gnd
rlabel metal1 4044 962 4296 978 0 _1560_.vdd
rlabel metal2 4193 813 4207 827 0 _1560_.D
rlabel metal2 4153 813 4167 827 0 _1560_.CLK
rlabel metal2 4073 813 4087 827 0 _1560_.Q
rlabel metal1 4284 722 4536 738 0 _1544_.gnd
rlabel metal1 4284 962 4536 978 0 _1544_.vdd
rlabel metal2 4373 813 4387 827 0 _1544_.D
rlabel metal2 4413 813 4427 827 0 _1544_.CLK
rlabel metal2 4493 813 4507 827 0 _1544_.Q
rlabel metal1 4524 722 4636 738 0 _850_.gnd
rlabel metal1 4524 962 4636 978 0 _850_.vdd
rlabel metal2 4533 813 4547 827 0 _850_.A
rlabel metal2 4553 833 4567 847 0 _850_.B
rlabel metal2 4593 833 4607 847 0 _850_.C
rlabel metal2 4573 813 4587 827 0 _850_.Y
rlabel nsubstratencontact 4756 968 4756 968 0 FILL71250x10950.vdd
rlabel metal1 4744 722 4776 738 0 FILL71250x10950.gnd
rlabel nsubstratencontact 4736 968 4736 968 0 FILL70950x10950.vdd
rlabel metal1 4724 722 4756 738 0 FILL70950x10950.gnd
rlabel metal1 4624 722 4736 738 0 _847_.gnd
rlabel metal1 4624 962 4736 978 0 _847_.vdd
rlabel metal2 4633 813 4647 827 0 _847_.A
rlabel metal2 4653 833 4667 847 0 _847_.B
rlabel metal2 4693 833 4707 847 0 _847_.C
rlabel metal2 4673 813 4687 827 0 _847_.Y
rlabel metal1 4 1202 116 1218 0 _1047_.gnd
rlabel metal1 4 962 116 978 0 _1047_.vdd
rlabel metal2 93 1113 107 1127 0 _1047_.A
rlabel metal2 73 1093 87 1107 0 _1047_.B
rlabel metal2 33 1093 47 1107 0 _1047_.C
rlabel metal2 53 1113 67 1127 0 _1047_.Y
rlabel metal1 104 1202 216 1218 0 _1043_.gnd
rlabel metal1 104 962 216 978 0 _1043_.vdd
rlabel metal2 113 1113 127 1127 0 _1043_.A
rlabel metal2 133 1093 147 1107 0 _1043_.B
rlabel metal2 173 1093 187 1107 0 _1043_.C
rlabel metal2 153 1113 167 1127 0 _1043_.Y
rlabel metal1 204 1202 316 1218 0 _1038_.gnd
rlabel metal1 204 962 316 978 0 _1038_.vdd
rlabel metal2 213 1093 227 1107 0 _1038_.A
rlabel metal2 233 1073 247 1087 0 _1038_.B
rlabel metal2 253 1093 267 1107 0 _1038_.C
rlabel metal2 273 1073 287 1087 0 _1038_.Y
rlabel metal1 304 1202 416 1218 0 _1075_.gnd
rlabel metal1 304 962 416 978 0 _1075_.vdd
rlabel metal2 313 1093 327 1107 0 _1075_.A
rlabel metal2 333 1133 347 1147 0 _1075_.B
rlabel metal2 353 1093 367 1107 0 _1075_.C
rlabel metal2 373 1113 387 1127 0 _1075_.Y
rlabel metal1 504 1202 616 1218 0 _1053_.gnd
rlabel metal1 504 962 616 978 0 _1053_.vdd
rlabel metal2 513 1093 527 1107 0 _1053_.A
rlabel metal2 533 1133 547 1147 0 _1053_.B
rlabel metal2 553 1093 567 1107 0 _1053_.C
rlabel metal2 573 1113 587 1127 0 _1053_.Y
rlabel metal1 404 1202 516 1218 0 _1044_.gnd
rlabel metal1 404 962 516 978 0 _1044_.vdd
rlabel metal2 413 1093 427 1107 0 _1044_.A
rlabel metal2 433 1073 447 1087 0 _1044_.B
rlabel metal2 453 1093 467 1107 0 _1044_.C
rlabel metal2 473 1073 487 1087 0 _1044_.Y
rlabel metal1 604 1202 696 1218 0 _1024_.gnd
rlabel metal1 604 962 696 978 0 _1024_.vdd
rlabel metal2 673 1073 687 1087 0 _1024_.A
rlabel metal2 633 1073 647 1087 0 _1024_.B
rlabel metal2 653 1093 667 1107 0 _1024_.Y
rlabel metal1 784 1202 896 1218 0 _1019_.gnd
rlabel metal1 784 962 896 978 0 _1019_.vdd
rlabel metal2 873 1093 887 1107 0 _1019_.A
rlabel metal2 853 1073 867 1087 0 _1019_.B
rlabel metal2 833 1093 847 1107 0 _1019_.C
rlabel metal2 813 1073 827 1087 0 _1019_.Y
rlabel metal1 684 1202 796 1218 0 _1045_.gnd
rlabel metal1 684 962 796 978 0 _1045_.vdd
rlabel metal2 773 1113 787 1127 0 _1045_.A
rlabel metal2 713 1113 727 1127 0 _1045_.Y
rlabel metal2 733 1073 747 1087 0 _1045_.B
rlabel metal1 984 1202 1096 1218 0 _1018_.gnd
rlabel metal1 984 962 1096 978 0 _1018_.vdd
rlabel metal2 993 1113 1007 1127 0 _1018_.A
rlabel metal2 1013 1093 1027 1107 0 _1018_.B
rlabel metal2 1053 1093 1067 1107 0 _1018_.C
rlabel metal2 1033 1113 1047 1127 0 _1018_.Y
rlabel metal1 884 1202 996 1218 0 _1016_.gnd
rlabel metal1 884 962 996 978 0 _1016_.vdd
rlabel metal2 973 1113 987 1127 0 _1016_.A
rlabel metal2 953 1093 967 1107 0 _1016_.B
rlabel metal2 913 1093 927 1107 0 _1016_.C
rlabel metal2 933 1113 947 1127 0 _1016_.Y
rlabel metal1 1084 1202 1196 1218 0 _961_.gnd
rlabel metal1 1084 962 1196 978 0 _961_.vdd
rlabel metal2 1173 1113 1187 1127 0 _961_.A
rlabel metal2 1153 1093 1167 1107 0 _961_.B
rlabel metal2 1113 1093 1127 1107 0 _961_.C
rlabel metal2 1133 1113 1147 1127 0 _961_.Y
rlabel metal1 1184 1202 1276 1218 0 _966_.gnd
rlabel metal1 1184 962 1276 978 0 _966_.vdd
rlabel metal2 1253 1073 1267 1087 0 _966_.A
rlabel metal2 1213 1073 1227 1087 0 _966_.B
rlabel metal2 1233 1093 1247 1107 0 _966_.Y
rlabel metal1 1264 1202 1376 1218 0 _960_.gnd
rlabel metal1 1264 962 1376 978 0 _960_.vdd
rlabel metal2 1353 1113 1367 1127 0 _960_.A
rlabel metal2 1293 1113 1307 1127 0 _960_.Y
rlabel metal2 1313 1073 1327 1087 0 _960_.B
rlabel metal1 1364 1202 1456 1218 0 _1014_.gnd
rlabel metal1 1364 962 1456 978 0 _1014_.vdd
rlabel metal2 1373 1073 1387 1087 0 _1014_.A
rlabel metal2 1413 1073 1427 1087 0 _1014_.B
rlabel metal2 1393 1093 1407 1107 0 _1014_.Y
rlabel metal1 1584 1202 1676 1218 0 _997_.gnd
rlabel metal1 1584 962 1676 978 0 _997_.vdd
rlabel metal2 1653 1073 1667 1087 0 _997_.A
rlabel metal2 1613 1073 1627 1087 0 _997_.B
rlabel metal2 1633 1093 1647 1107 0 _997_.Y
rlabel metal1 1504 1202 1596 1218 0 _993_.gnd
rlabel metal1 1504 962 1596 978 0 _993_.vdd
rlabel metal2 1573 1073 1587 1087 0 _993_.A
rlabel metal2 1533 1073 1547 1087 0 _993_.B
rlabel metal2 1553 1093 1567 1107 0 _993_.Y
rlabel metal1 1444 1202 1516 1218 0 _934_.gnd
rlabel metal1 1444 962 1516 978 0 _934_.vdd
rlabel metal2 1493 1093 1507 1107 0 _934_.A
rlabel metal2 1473 1113 1487 1127 0 _934_.Y
rlabel metal1 1764 1202 1856 1218 0 _994_.gnd
rlabel metal1 1764 962 1856 978 0 _994_.vdd
rlabel metal2 1833 1073 1847 1087 0 _994_.A
rlabel metal2 1793 1073 1807 1087 0 _994_.B
rlabel metal2 1813 1093 1827 1107 0 _994_.Y
rlabel metal1 1844 1202 1956 1218 0 _995_.gnd
rlabel metal1 1844 962 1956 978 0 _995_.vdd
rlabel metal2 1853 1093 1867 1107 0 _995_.A
rlabel metal2 1873 1073 1887 1087 0 _995_.B
rlabel metal2 1893 1093 1907 1107 0 _995_.C
rlabel metal2 1913 1073 1927 1087 0 _995_.Y
rlabel metal1 1664 1202 1776 1218 0 _991_.gnd
rlabel metal1 1664 962 1776 978 0 _991_.vdd
rlabel metal2 1673 1093 1687 1107 0 _991_.A
rlabel metal2 1693 1073 1707 1087 0 _991_.B
rlabel metal2 1713 1093 1727 1107 0 _991_.C
rlabel metal2 1733 1073 1747 1087 0 _991_.Y
rlabel metal1 1944 1202 2036 1218 0 _955_.gnd
rlabel metal1 1944 962 2036 978 0 _955_.vdd
rlabel metal2 1953 1073 1967 1087 0 _955_.A
rlabel metal2 1993 1073 2007 1087 0 _955_.B
rlabel metal2 1973 1093 1987 1107 0 _955_.Y
rlabel metal1 2024 1202 2156 1218 0 _1002_.gnd
rlabel metal1 2024 962 2156 978 0 _1002_.vdd
rlabel metal2 2133 1113 2147 1127 0 _1002_.A
rlabel metal2 2113 1093 2127 1107 0 _1002_.B
rlabel metal2 2053 1113 2067 1127 0 _1002_.C
rlabel metal2 2073 1093 2087 1107 0 _1002_.D
rlabel metal2 2093 1113 2107 1127 0 _1002_.Y
rlabel metal1 2244 1202 2336 1218 0 _1000_.gnd
rlabel metal1 2244 962 2336 978 0 _1000_.vdd
rlabel metal2 2313 1073 2327 1087 0 _1000_.A
rlabel metal2 2273 1073 2287 1087 0 _1000_.B
rlabel metal2 2293 1093 2307 1107 0 _1000_.Y
rlabel metal1 2324 1202 2436 1218 0 _949_.gnd
rlabel metal1 2324 962 2436 978 0 _949_.vdd
rlabel metal2 2333 1093 2347 1107 0 _949_.A
rlabel metal2 2353 1133 2367 1147 0 _949_.B
rlabel metal2 2373 1093 2387 1107 0 _949_.C
rlabel metal2 2393 1113 2407 1127 0 _949_.Y
rlabel metal1 2144 1202 2256 1218 0 _950_.gnd
rlabel metal1 2144 962 2256 978 0 _950_.vdd
rlabel metal2 2233 1093 2247 1107 0 _950_.A
rlabel metal2 2213 1073 2227 1087 0 _950_.B
rlabel metal2 2193 1093 2207 1107 0 _950_.C
rlabel metal2 2173 1073 2187 1087 0 _950_.Y
rlabel metal1 2484 1202 2576 1218 0 _951_.gnd
rlabel metal1 2484 962 2576 978 0 _951_.vdd
rlabel metal2 2553 1073 2567 1087 0 _951_.A
rlabel metal2 2513 1073 2527 1087 0 _951_.B
rlabel metal2 2533 1093 2547 1107 0 _951_.Y
rlabel metal1 2424 1202 2496 1218 0 _914_.gnd
rlabel metal1 2424 962 2496 978 0 _914_.vdd
rlabel metal2 2473 1133 2487 1147 0 _914_.A
rlabel metal2 2453 1093 2467 1107 0 _914_.Y
rlabel metal1 2564 1202 2696 1218 0 _952_.gnd
rlabel metal1 2564 962 2696 978 0 _952_.vdd
rlabel metal2 2673 1113 2687 1127 0 _952_.A
rlabel metal2 2653 1093 2667 1107 0 _952_.B
rlabel metal2 2593 1113 2607 1127 0 _952_.C
rlabel metal2 2633 1113 2647 1127 0 _952_.Y
rlabel metal2 2613 1093 2627 1107 0 _952_.D
rlabel metal1 2684 1202 2776 1218 0 BUFX2_insert0.gnd
rlabel metal1 2684 962 2776 978 0 BUFX2_insert0.vdd
rlabel metal2 2693 1113 2707 1127 0 BUFX2_insert0.A
rlabel metal2 2733 1113 2747 1127 0 BUFX2_insert0.Y
rlabel metal1 2764 1202 3016 1218 0 _1550_.gnd
rlabel metal1 2764 962 3016 978 0 _1550_.vdd
rlabel metal2 2853 1113 2867 1127 0 _1550_.D
rlabel metal2 2893 1113 2907 1127 0 _1550_.CLK
rlabel metal2 2973 1113 2987 1127 0 _1550_.Q
rlabel metal1 3084 1202 3196 1218 0 _814_.gnd
rlabel metal1 3084 962 3196 978 0 _814_.vdd
rlabel metal2 3173 1113 3187 1127 0 _814_.A
rlabel metal2 3153 1093 3167 1107 0 _814_.B
rlabel metal2 3113 1093 3127 1107 0 _814_.C
rlabel metal2 3133 1113 3147 1127 0 _814_.Y
rlabel metal1 3004 1202 3096 1218 0 _813_.gnd
rlabel metal1 3004 962 3096 978 0 _813_.vdd
rlabel metal2 3013 1073 3027 1087 0 _813_.A
rlabel metal2 3053 1073 3067 1087 0 _813_.B
rlabel metal2 3033 1093 3047 1107 0 _813_.Y
rlabel metal1 3184 1202 3316 1218 0 _1197_.gnd
rlabel metal1 3184 962 3316 978 0 _1197_.vdd
rlabel metal2 3213 1113 3227 1127 0 _1197_.A
rlabel metal2 3253 1113 3267 1127 0 _1197_.Y
rlabel metal1 3464 1202 3676 1218 0 CLKBUF1_insert15.gnd
rlabel metal1 3464 962 3676 978 0 CLKBUF1_insert15.vdd
rlabel metal2 3493 1093 3507 1107 0 CLKBUF1_insert15.A
rlabel metal2 3633 1093 3647 1107 0 CLKBUF1_insert15.Y
rlabel metal1 3384 1202 3476 1218 0 BUFX2_insert4.gnd
rlabel metal1 3384 962 3476 978 0 BUFX2_insert4.vdd
rlabel metal2 3393 1113 3407 1127 0 BUFX2_insert4.A
rlabel metal2 3433 1113 3447 1127 0 BUFX2_insert4.Y
rlabel metal1 3304 1202 3396 1218 0 BUFX2_insert2.gnd
rlabel metal1 3304 962 3396 978 0 BUFX2_insert2.vdd
rlabel metal2 3373 1113 3387 1127 0 BUFX2_insert2.A
rlabel metal2 3333 1113 3347 1127 0 BUFX2_insert2.Y
rlabel metal1 3664 1202 3876 1218 0 CLKBUF1_insert13.gnd
rlabel metal1 3664 962 3876 978 0 CLKBUF1_insert13.vdd
rlabel metal2 3693 1093 3707 1107 0 CLKBUF1_insert13.A
rlabel metal2 3833 1093 3847 1107 0 CLKBUF1_insert13.Y
rlabel metal1 3864 1202 3956 1218 0 BUFX2_insert20.gnd
rlabel metal1 3864 962 3956 978 0 BUFX2_insert20.vdd
rlabel metal2 3873 1113 3887 1127 0 BUFX2_insert20.A
rlabel metal2 3913 1113 3927 1127 0 BUFX2_insert20.Y
rlabel metal1 3944 1202 4036 1218 0 _1330_.gnd
rlabel metal1 3944 962 4036 978 0 _1330_.vdd
rlabel metal2 3953 1073 3967 1087 0 _1330_.A
rlabel metal2 3993 1073 4007 1087 0 _1330_.B
rlabel metal2 3973 1093 3987 1107 0 _1330_.Y
rlabel metal1 4024 1202 4276 1218 0 _1575_.gnd
rlabel metal1 4024 962 4276 978 0 _1575_.vdd
rlabel metal2 4173 1113 4187 1127 0 _1575_.D
rlabel metal2 4133 1113 4147 1127 0 _1575_.CLK
rlabel metal2 4053 1113 4067 1127 0 _1575_.Q
rlabel metal1 4264 1202 4356 1218 0 _1474_.gnd
rlabel metal1 4264 962 4356 978 0 _1474_.vdd
rlabel metal2 4273 1073 4287 1087 0 _1474_.A
rlabel metal2 4313 1073 4327 1087 0 _1474_.B
rlabel metal2 4293 1093 4307 1107 0 _1474_.Y
rlabel metal1 4344 1202 4456 1218 0 _1478_.gnd
rlabel metal1 4344 962 4456 978 0 _1478_.vdd
rlabel metal2 4353 1113 4367 1127 0 _1478_.A
rlabel metal2 4373 1093 4387 1107 0 _1478_.B
rlabel metal2 4413 1093 4427 1107 0 _1478_.C
rlabel metal2 4393 1113 4407 1127 0 _1478_.Y
rlabel metal1 4524 1202 4636 1218 0 _1476_.gnd
rlabel metal1 4524 962 4636 978 0 _1476_.vdd
rlabel metal2 4533 1113 4547 1127 0 _1476_.A
rlabel metal2 4553 1093 4567 1107 0 _1476_.B
rlabel metal2 4593 1093 4607 1107 0 _1476_.C
rlabel metal2 4573 1113 4587 1127 0 _1476_.Y
rlabel metal1 4444 1202 4536 1218 0 _1477_.gnd
rlabel metal1 4444 962 4536 978 0 _1477_.vdd
rlabel metal2 4513 1073 4527 1087 0 _1477_.A
rlabel metal2 4473 1073 4487 1087 0 _1477_.B
rlabel metal2 4493 1093 4507 1107 0 _1477_.Y
rlabel nsubstratencontact 4764 972 4764 972 0 FILL71250x14550.vdd
rlabel metal1 4744 1202 4776 1218 0 FILL71250x14550.gnd
rlabel nsubstratencontact 4744 972 4744 972 0 FILL70950x14550.vdd
rlabel metal1 4724 1202 4756 1218 0 FILL70950x14550.gnd
rlabel metal1 4624 1202 4736 1218 0 _1475_.gnd
rlabel metal1 4624 962 4736 978 0 _1475_.vdd
rlabel metal2 4633 1093 4647 1107 0 _1475_.A
rlabel metal2 4653 1073 4667 1087 0 _1475_.B
rlabel metal2 4673 1093 4687 1107 0 _1475_.C
rlabel metal2 4693 1073 4707 1087 0 _1475_.Y
rlabel metal1 4 1202 116 1218 0 _1042_.gnd
rlabel metal1 4 1442 116 1458 0 _1042_.vdd
rlabel metal2 93 1313 107 1327 0 _1042_.A
rlabel metal2 73 1273 87 1287 0 _1042_.B
rlabel metal2 53 1313 67 1327 0 _1042_.C
rlabel metal2 33 1293 47 1307 0 _1042_.Y
rlabel metal1 204 1202 316 1218 0 _1046_.gnd
rlabel metal1 204 1442 316 1458 0 _1046_.vdd
rlabel metal2 213 1313 227 1327 0 _1046_.A
rlabel metal2 233 1333 247 1347 0 _1046_.B
rlabel metal2 253 1313 267 1327 0 _1046_.C
rlabel metal2 273 1333 287 1347 0 _1046_.Y
rlabel metal1 104 1202 216 1218 0 _1032_.gnd
rlabel metal1 104 1442 216 1458 0 _1032_.vdd
rlabel metal2 113 1313 127 1327 0 _1032_.A
rlabel metal2 133 1333 147 1347 0 _1032_.B
rlabel metal2 153 1313 167 1327 0 _1032_.C
rlabel metal2 173 1333 187 1347 0 _1032_.Y
rlabel metal1 384 1202 496 1218 0 _1076_.gnd
rlabel metal1 384 1442 496 1458 0 _1076_.vdd
rlabel metal2 393 1293 407 1307 0 _1076_.A
rlabel metal2 413 1313 427 1327 0 _1076_.B
rlabel metal2 453 1313 467 1327 0 _1076_.C
rlabel metal2 433 1293 447 1307 0 _1076_.Y
rlabel metal1 304 1202 396 1218 0 _1027_.gnd
rlabel metal1 304 1442 396 1458 0 _1027_.vdd
rlabel metal2 373 1333 387 1347 0 _1027_.A
rlabel metal2 333 1333 347 1347 0 _1027_.B
rlabel metal2 353 1313 367 1327 0 _1027_.Y
rlabel metal1 484 1202 596 1218 0 _1052_.gnd
rlabel metal1 484 1442 596 1458 0 _1052_.vdd
rlabel metal2 493 1313 507 1327 0 _1052_.A
rlabel metal2 513 1273 527 1287 0 _1052_.B
rlabel metal2 533 1313 547 1327 0 _1052_.C
rlabel metal2 553 1293 567 1307 0 _1052_.Y
rlabel metal1 584 1202 696 1218 0 _1057_.gnd
rlabel metal1 584 1442 696 1458 0 _1057_.vdd
rlabel metal2 593 1293 607 1307 0 _1057_.A
rlabel metal2 613 1313 627 1327 0 _1057_.B
rlabel metal2 653 1313 667 1327 0 _1057_.C
rlabel metal2 633 1293 647 1307 0 _1057_.Y
rlabel metal1 684 1202 796 1218 0 _1054_.gnd
rlabel metal1 684 1442 796 1458 0 _1054_.vdd
rlabel metal2 693 1293 707 1307 0 _1054_.A
rlabel metal2 713 1313 727 1327 0 _1054_.B
rlabel metal2 753 1313 767 1327 0 _1054_.C
rlabel metal2 733 1293 747 1307 0 _1054_.Y
rlabel metal1 784 1202 896 1218 0 _1015_.gnd
rlabel metal1 784 1442 896 1458 0 _1015_.vdd
rlabel metal2 793 1293 807 1307 0 _1015_.A
rlabel metal2 853 1293 867 1307 0 _1015_.Y
rlabel metal2 833 1333 847 1347 0 _1015_.B
rlabel metal1 964 1202 1056 1218 0 _1074_.gnd
rlabel metal1 964 1442 1056 1458 0 _1074_.vdd
rlabel metal2 973 1333 987 1347 0 _1074_.A
rlabel metal2 1013 1333 1027 1347 0 _1074_.B
rlabel metal2 993 1313 1007 1327 0 _1074_.Y
rlabel metal1 884 1202 976 1218 0 _1021_.gnd
rlabel metal1 884 1442 976 1458 0 _1021_.vdd
rlabel metal2 953 1333 967 1347 0 _1021_.A
rlabel metal2 913 1333 927 1347 0 _1021_.B
rlabel metal2 933 1313 947 1327 0 _1021_.Y
rlabel metal1 1044 1202 1156 1218 0 _1023_.gnd
rlabel metal1 1044 1442 1156 1458 0 _1023_.vdd
rlabel metal2 1133 1313 1147 1327 0 _1023_.A
rlabel metal2 1113 1333 1127 1347 0 _1023_.B
rlabel metal2 1093 1313 1107 1327 0 _1023_.C
rlabel metal2 1073 1333 1087 1347 0 _1023_.Y
rlabel metal1 1304 1202 1416 1218 0 _1022_.gnd
rlabel metal1 1304 1442 1416 1458 0 _1022_.vdd
rlabel metal2 1313 1293 1327 1307 0 _1022_.A
rlabel metal2 1333 1313 1347 1327 0 _1022_.B
rlabel metal2 1373 1313 1387 1327 0 _1022_.C
rlabel metal2 1353 1293 1367 1307 0 _1022_.Y
rlabel metal1 1144 1202 1216 1218 0 _1020_.gnd
rlabel metal1 1144 1442 1216 1458 0 _1020_.vdd
rlabel metal2 1193 1273 1207 1287 0 _1020_.A
rlabel metal2 1173 1313 1187 1327 0 _1020_.Y
rlabel metal1 1204 1202 1316 1218 0 _1017_.gnd
rlabel metal1 1204 1442 1316 1458 0 _1017_.vdd
rlabel metal2 1293 1293 1307 1307 0 _1017_.A
rlabel metal2 1233 1293 1247 1307 0 _1017_.Y
rlabel metal2 1253 1333 1267 1347 0 _1017_.B
rlabel metal1 1404 1202 1516 1218 0 _1010_.gnd
rlabel metal1 1404 1442 1516 1458 0 _1010_.vdd
rlabel metal2 1493 1293 1507 1307 0 _1010_.A
rlabel metal2 1473 1313 1487 1327 0 _1010_.B
rlabel metal2 1433 1313 1447 1327 0 _1010_.C
rlabel metal2 1453 1293 1467 1307 0 _1010_.Y
rlabel metal1 1584 1202 1696 1218 0 _936_.gnd
rlabel metal1 1584 1442 1696 1458 0 _936_.vdd
rlabel metal2 1593 1293 1607 1307 0 _936_.A
rlabel metal2 1613 1313 1627 1327 0 _936_.B
rlabel metal2 1653 1313 1667 1327 0 _936_.C
rlabel metal2 1633 1293 1647 1307 0 _936_.Y
rlabel metal1 1504 1202 1596 1218 0 _1009_.gnd
rlabel metal1 1504 1442 1596 1458 0 _1009_.vdd
rlabel metal2 1513 1333 1527 1347 0 _1009_.A
rlabel metal2 1553 1333 1567 1347 0 _1009_.B
rlabel metal2 1533 1313 1547 1327 0 _1009_.Y
rlabel metal1 1684 1202 1776 1218 0 _935_.gnd
rlabel metal1 1684 1442 1776 1458 0 _935_.vdd
rlabel metal2 1693 1333 1707 1347 0 _935_.A
rlabel metal2 1733 1333 1747 1347 0 _935_.B
rlabel metal2 1713 1313 1727 1327 0 _935_.Y
rlabel metal1 1764 1202 1876 1218 0 _1007_.gnd
rlabel metal1 1764 1442 1876 1458 0 _1007_.vdd
rlabel metal2 1773 1313 1787 1327 0 _1007_.A
rlabel metal2 1793 1273 1807 1287 0 _1007_.B
rlabel metal2 1813 1313 1827 1327 0 _1007_.C
rlabel metal2 1833 1293 1847 1307 0 _1007_.Y
rlabel metal1 1864 1202 1976 1218 0 _996_.gnd
rlabel metal1 1864 1442 1976 1458 0 _996_.vdd
rlabel metal2 1873 1313 1887 1327 0 _996_.A
rlabel metal2 1893 1333 1907 1347 0 _996_.B
rlabel metal2 1913 1313 1927 1327 0 _996_.C
rlabel metal2 1933 1333 1947 1347 0 _996_.Y
rlabel metal1 1964 1202 2076 1218 0 _1008_.gnd
rlabel metal1 1964 1442 2076 1458 0 _1008_.vdd
rlabel metal2 1973 1293 1987 1307 0 _1008_.A
rlabel metal2 1993 1313 2007 1327 0 _1008_.B
rlabel metal2 2033 1313 2047 1327 0 _1008_.C
rlabel metal2 2013 1293 2027 1307 0 _1008_.Y
rlabel metal1 2064 1202 2136 1218 0 _956_.gnd
rlabel metal1 2064 1442 2136 1458 0 _956_.vdd
rlabel metal2 2073 1273 2087 1287 0 _956_.A
rlabel metal2 2093 1313 2107 1327 0 _956_.Y
rlabel metal1 2124 1202 2236 1218 0 _998_.gnd
rlabel metal1 2124 1442 2236 1458 0 _998_.vdd
rlabel metal2 2133 1313 2147 1327 0 _998_.A
rlabel metal2 2153 1333 2167 1347 0 _998_.B
rlabel metal2 2173 1313 2187 1327 0 _998_.C
rlabel metal2 2193 1333 2207 1347 0 _998_.Y
rlabel metal1 2404 1202 2496 1218 0 _1308_.gnd
rlabel metal1 2404 1442 2496 1458 0 _1308_.vdd
rlabel metal2 2473 1333 2487 1347 0 _1308_.A
rlabel metal2 2433 1333 2447 1347 0 _1308_.B
rlabel metal2 2453 1313 2467 1327 0 _1308_.Y
rlabel metal1 2224 1202 2316 1218 0 _999_.gnd
rlabel metal1 2224 1442 2316 1458 0 _999_.vdd
rlabel metal2 2233 1333 2247 1347 0 _999_.A
rlabel metal2 2273 1333 2287 1347 0 _999_.B
rlabel metal2 2253 1313 2267 1327 0 _999_.Y
rlabel metal1 2304 1202 2416 1218 0 _1001_.gnd
rlabel metal1 2304 1442 2416 1458 0 _1001_.vdd
rlabel metal2 2313 1273 2327 1287 0 _1001_.A
rlabel metal2 2333 1293 2347 1307 0 _1001_.B
rlabel metal2 2373 1313 2387 1327 0 _1001_.Y
rlabel metal1 2544 1202 2636 1218 0 BUFX2_insert7.gnd
rlabel metal1 2544 1442 2636 1458 0 BUFX2_insert7.vdd
rlabel metal2 2613 1293 2627 1307 0 BUFX2_insert7.A
rlabel metal2 2573 1293 2587 1307 0 BUFX2_insert7.Y
rlabel metal1 2624 1202 2736 1218 0 _1310_.gnd
rlabel metal1 2624 1442 2736 1458 0 _1310_.vdd
rlabel metal2 2633 1293 2647 1307 0 _1310_.A
rlabel metal2 2653 1313 2667 1327 0 _1310_.B
rlabel metal2 2693 1313 2707 1327 0 _1310_.C
rlabel metal2 2673 1293 2687 1307 0 _1310_.Y
rlabel metal1 2484 1202 2556 1218 0 _1309_.gnd
rlabel metal1 2484 1442 2556 1458 0 _1309_.vdd
rlabel metal2 2493 1273 2507 1287 0 _1309_.A
rlabel metal2 2513 1313 2527 1327 0 _1309_.Y
rlabel metal1 2844 1202 3096 1218 0 _1591_.gnd
rlabel metal1 2844 1442 3096 1458 0 _1591_.vdd
rlabel metal2 2933 1293 2947 1307 0 _1591_.D
rlabel metal2 2973 1293 2987 1307 0 _1591_.CLK
rlabel metal2 3053 1293 3067 1307 0 _1591_.Q
rlabel metal1 2724 1202 2856 1218 0 _1311_.gnd
rlabel metal1 2724 1442 2856 1458 0 _1311_.vdd
rlabel metal2 2833 1293 2847 1307 0 _1311_.A
rlabel metal2 2813 1313 2827 1327 0 _1311_.B
rlabel metal2 2753 1293 2767 1307 0 _1311_.C
rlabel metal2 2793 1293 2807 1307 0 _1311_.Y
rlabel metal2 2773 1313 2787 1327 0 _1311_.D
rlabel metal1 3164 1202 3276 1218 0 _1517_.gnd
rlabel metal1 3164 1442 3276 1458 0 _1517_.vdd
rlabel metal2 3253 1313 3267 1327 0 _1517_.A
rlabel metal2 3233 1273 3247 1287 0 _1517_.B
rlabel metal2 3213 1313 3227 1327 0 _1517_.C
rlabel metal2 3193 1293 3207 1307 0 _1517_.Y
rlabel metal1 3084 1202 3176 1218 0 _1516_.gnd
rlabel metal1 3084 1442 3176 1458 0 _1516_.vdd
rlabel metal2 3113 1293 3127 1307 0 _1516_.B
rlabel metal2 3153 1293 3167 1307 0 _1516_.A
rlabel metal2 3133 1273 3147 1287 0 _1516_.Y
rlabel metal1 3264 1202 3516 1218 0 _1558_.gnd
rlabel metal1 3264 1442 3516 1458 0 _1558_.vdd
rlabel metal2 3353 1293 3367 1307 0 _1558_.D
rlabel metal2 3393 1293 3407 1307 0 _1558_.CLK
rlabel metal2 3473 1293 3487 1307 0 _1558_.Q
rlabel metal1 3564 1202 3656 1218 0 _1447_.gnd
rlabel metal1 3564 1442 3656 1458 0 _1447_.vdd
rlabel metal2 3593 1293 3607 1307 0 _1447_.B
rlabel metal2 3633 1293 3647 1307 0 _1447_.A
rlabel metal2 3613 1273 3627 1287 0 _1447_.Y
rlabel metal1 3644 1202 3736 1218 0 _1446_.gnd
rlabel metal1 3644 1442 3736 1458 0 _1446_.vdd
rlabel metal2 3673 1293 3687 1307 0 _1446_.B
rlabel metal2 3713 1293 3727 1307 0 _1446_.A
rlabel metal2 3693 1273 3707 1287 0 _1446_.Y
rlabel metal1 3504 1202 3576 1218 0 _1295_.gnd
rlabel metal1 3504 1442 3576 1458 0 _1295_.vdd
rlabel metal2 3553 1273 3567 1287 0 _1295_.A
rlabel metal2 3533 1313 3547 1327 0 _1295_.Y
rlabel metal1 3724 1202 3796 1218 0 _839_.gnd
rlabel metal1 3724 1442 3796 1458 0 _839_.vdd
rlabel metal2 3733 1273 3747 1287 0 _839_.A
rlabel metal2 3753 1313 3767 1327 0 _839_.Y
rlabel metal1 3784 1202 4036 1218 0 _1542_.gnd
rlabel metal1 3784 1442 4036 1458 0 _1542_.vdd
rlabel metal2 3933 1293 3947 1307 0 _1542_.D
rlabel metal2 3893 1293 3907 1307 0 _1542_.CLK
rlabel metal2 3813 1293 3827 1307 0 _1542_.Q
rlabel metal1 4204 1202 4296 1218 0 BUFX2_insert6.gnd
rlabel metal1 4204 1442 4296 1458 0 BUFX2_insert6.vdd
rlabel metal2 4273 1293 4287 1307 0 BUFX2_insert6.A
rlabel metal2 4233 1293 4247 1307 0 BUFX2_insert6.Y
rlabel metal1 4024 1202 4136 1218 0 _841_.gnd
rlabel metal1 4024 1442 4136 1458 0 _841_.vdd
rlabel metal2 4033 1293 4047 1307 0 _841_.A
rlabel metal2 4053 1313 4067 1327 0 _841_.B
rlabel metal2 4093 1313 4107 1327 0 _841_.C
rlabel metal2 4073 1293 4087 1307 0 _841_.Y
rlabel metal1 4124 1202 4216 1218 0 _840_.gnd
rlabel metal1 4124 1442 4216 1458 0 _840_.vdd
rlabel metal2 4133 1333 4147 1347 0 _840_.A
rlabel metal2 4173 1333 4187 1347 0 _840_.B
rlabel metal2 4153 1313 4167 1327 0 _840_.Y
rlabel metal1 4364 1202 4476 1218 0 _1473_.gnd
rlabel metal1 4364 1442 4476 1458 0 _1473_.vdd
rlabel metal2 4453 1293 4467 1307 0 _1473_.A
rlabel metal2 4433 1313 4447 1327 0 _1473_.B
rlabel metal2 4393 1313 4407 1327 0 _1473_.C
rlabel metal2 4413 1293 4427 1307 0 _1473_.Y
rlabel metal1 4464 1202 4576 1218 0 _1472_.gnd
rlabel metal1 4464 1442 4576 1458 0 _1472_.vdd
rlabel metal2 4553 1293 4567 1307 0 _1472_.A
rlabel metal2 4533 1313 4547 1327 0 _1472_.B
rlabel metal2 4493 1313 4507 1327 0 _1472_.C
rlabel metal2 4513 1293 4527 1307 0 _1472_.Y
rlabel metal1 4284 1202 4376 1218 0 _1464_.gnd
rlabel metal1 4284 1442 4376 1458 0 _1464_.vdd
rlabel metal2 4353 1333 4367 1347 0 _1464_.A
rlabel metal2 4313 1333 4327 1347 0 _1464_.B
rlabel metal2 4333 1313 4347 1327 0 _1464_.Y
rlabel metal1 4564 1202 4656 1218 0 _1469_.gnd
rlabel metal1 4564 1442 4656 1458 0 _1469_.vdd
rlabel metal2 4613 1293 4627 1307 0 _1469_.B
rlabel metal2 4573 1293 4587 1307 0 _1469_.A
rlabel metal2 4593 1273 4607 1287 0 _1469_.Y
rlabel metal1 4704 1202 4776 1218 0 _1489_.gnd
rlabel metal1 4704 1442 4776 1458 0 _1489_.vdd
rlabel metal2 4753 1273 4767 1287 0 _1489_.A
rlabel metal2 4733 1313 4747 1327 0 _1489_.Y
rlabel metal1 4644 1202 4716 1218 0 _845_.gnd
rlabel metal1 4644 1442 4716 1458 0 _845_.vdd
rlabel metal2 4653 1273 4667 1287 0 _845_.A
rlabel metal2 4673 1313 4687 1327 0 _845_.Y
rlabel metal1 264 1682 356 1698 0 _1035_.gnd
rlabel metal1 264 1442 356 1458 0 _1035_.vdd
rlabel metal2 273 1553 287 1567 0 _1035_.A
rlabel metal2 313 1553 327 1567 0 _1035_.B
rlabel metal2 293 1573 307 1587 0 _1035_.Y
rlabel metal1 64 1682 176 1698 0 _1041_.gnd
rlabel metal1 64 1442 176 1458 0 _1041_.vdd
rlabel metal2 153 1573 167 1587 0 _1041_.A
rlabel metal2 133 1613 147 1627 0 _1041_.B
rlabel metal2 113 1573 127 1587 0 _1041_.C
rlabel metal2 93 1593 107 1607 0 _1041_.Y
rlabel metal1 4 1682 76 1698 0 _1033_.gnd
rlabel metal1 4 1442 76 1458 0 _1033_.vdd
rlabel metal2 53 1613 67 1627 0 _1033_.A
rlabel metal2 33 1573 47 1587 0 _1033_.Y
rlabel metal1 164 1682 276 1698 0 _1037_.gnd
rlabel metal1 164 1442 276 1458 0 _1037_.vdd
rlabel metal2 173 1573 187 1587 0 _1037_.A
rlabel metal2 193 1553 207 1567 0 _1037_.B
rlabel metal2 213 1573 227 1587 0 _1037_.C
rlabel metal2 233 1553 247 1567 0 _1037_.Y
rlabel metal1 444 1682 536 1698 0 BUFX2_insert21.gnd
rlabel metal1 444 1442 536 1458 0 BUFX2_insert21.vdd
rlabel metal2 513 1593 527 1607 0 BUFX2_insert21.A
rlabel metal2 473 1593 487 1607 0 BUFX2_insert21.Y
rlabel metal1 344 1682 456 1698 0 _1102_.gnd
rlabel metal1 344 1442 456 1458 0 _1102_.vdd
rlabel metal2 433 1593 447 1607 0 _1102_.A
rlabel metal2 413 1573 427 1587 0 _1102_.B
rlabel metal2 373 1573 387 1587 0 _1102_.C
rlabel metal2 393 1593 407 1607 0 _1102_.Y
rlabel metal1 524 1682 596 1698 0 _1112_.gnd
rlabel metal1 524 1442 596 1458 0 _1112_.vdd
rlabel metal2 573 1613 587 1627 0 _1112_.A
rlabel metal2 553 1573 567 1587 0 _1112_.Y
rlabel metal1 684 1682 796 1698 0 _1113_.gnd
rlabel metal1 684 1442 796 1458 0 _1113_.vdd
rlabel metal2 693 1573 707 1587 0 _1113_.A
rlabel metal2 713 1613 727 1627 0 _1113_.B
rlabel metal2 733 1573 747 1587 0 _1113_.C
rlabel metal2 753 1593 767 1607 0 _1113_.Y
rlabel metal1 784 1682 896 1698 0 _1049_.gnd
rlabel metal1 784 1442 896 1458 0 _1049_.vdd
rlabel metal2 793 1573 807 1587 0 _1049_.A
rlabel metal2 813 1553 827 1567 0 _1049_.B
rlabel metal2 833 1573 847 1587 0 _1049_.C
rlabel metal2 853 1553 867 1567 0 _1049_.Y
rlabel metal1 584 1682 696 1698 0 _1048_.gnd
rlabel metal1 584 1442 696 1458 0 _1048_.vdd
rlabel metal2 593 1573 607 1587 0 _1048_.A
rlabel metal2 613 1553 627 1567 0 _1048_.B
rlabel metal2 633 1573 647 1587 0 _1048_.C
rlabel metal2 653 1553 667 1567 0 _1048_.Y
rlabel metal1 884 1682 996 1698 0 _1072_.gnd
rlabel metal1 884 1442 996 1458 0 _1072_.vdd
rlabel metal2 893 1573 907 1587 0 _1072_.A
rlabel metal2 913 1613 927 1627 0 _1072_.B
rlabel metal2 933 1573 947 1587 0 _1072_.C
rlabel metal2 953 1593 967 1607 0 _1072_.Y
rlabel metal1 984 1682 1096 1698 0 _1056_.gnd
rlabel metal1 984 1442 1096 1458 0 _1056_.vdd
rlabel metal2 993 1573 1007 1587 0 _1056_.A
rlabel metal2 1013 1553 1027 1567 0 _1056_.B
rlabel metal2 1033 1573 1047 1587 0 _1056_.C
rlabel metal2 1053 1553 1067 1567 0 _1056_.Y
rlabel metal1 1084 1682 1196 1698 0 _1073_.gnd
rlabel metal1 1084 1442 1196 1458 0 _1073_.vdd
rlabel metal2 1173 1593 1187 1607 0 _1073_.A
rlabel metal2 1153 1573 1167 1587 0 _1073_.B
rlabel metal2 1113 1573 1127 1587 0 _1073_.C
rlabel metal2 1133 1593 1147 1607 0 _1073_.Y
rlabel metal1 1284 1682 1396 1698 0 _1063_.gnd
rlabel metal1 1284 1442 1396 1458 0 _1063_.vdd
rlabel metal2 1293 1573 1307 1587 0 _1063_.A
rlabel metal2 1313 1613 1327 1627 0 _1063_.B
rlabel metal2 1333 1573 1347 1587 0 _1063_.C
rlabel metal2 1353 1593 1367 1607 0 _1063_.Y
rlabel metal1 1184 1682 1296 1698 0 _1055_.gnd
rlabel metal1 1184 1442 1296 1458 0 _1055_.vdd
rlabel metal2 1193 1573 1207 1587 0 _1055_.A
rlabel metal2 1213 1553 1227 1567 0 _1055_.B
rlabel metal2 1233 1573 1247 1587 0 _1055_.C
rlabel metal2 1253 1553 1267 1567 0 _1055_.Y
rlabel metal1 1544 1682 1656 1698 0 _1062_.gnd
rlabel metal1 1544 1442 1656 1458 0 _1062_.vdd
rlabel metal2 1553 1573 1567 1587 0 _1062_.A
rlabel metal2 1573 1613 1587 1627 0 _1062_.B
rlabel metal2 1593 1573 1607 1587 0 _1062_.C
rlabel metal2 1613 1593 1627 1607 0 _1062_.Y
rlabel metal1 1384 1682 1456 1698 0 _1011_.gnd
rlabel metal1 1384 1442 1456 1458 0 _1011_.vdd
rlabel metal2 1433 1613 1447 1627 0 _1011_.A
rlabel metal2 1413 1573 1427 1587 0 _1011_.Y
rlabel metal1 1444 1682 1556 1698 0 _1058_.gnd
rlabel metal1 1444 1442 1556 1458 0 _1058_.vdd
rlabel metal2 1453 1573 1467 1587 0 _1058_.A
rlabel metal2 1473 1553 1487 1567 0 _1058_.B
rlabel metal2 1493 1573 1507 1587 0 _1058_.C
rlabel metal2 1513 1553 1527 1567 0 _1058_.Y
rlabel metal1 1744 1682 1856 1698 0 _1064_.gnd
rlabel metal1 1744 1442 1856 1458 0 _1064_.vdd
rlabel metal2 1753 1593 1767 1607 0 _1064_.A
rlabel metal2 1773 1573 1787 1587 0 _1064_.B
rlabel metal2 1813 1573 1827 1587 0 _1064_.C
rlabel metal2 1793 1593 1807 1607 0 _1064_.Y
rlabel metal1 1844 1682 1956 1698 0 _1061_.gnd
rlabel metal1 1844 1442 1956 1458 0 _1061_.vdd
rlabel metal2 1933 1573 1947 1587 0 _1061_.A
rlabel metal2 1913 1613 1927 1627 0 _1061_.B
rlabel metal2 1893 1573 1907 1587 0 _1061_.C
rlabel metal2 1873 1593 1887 1607 0 _1061_.Y
rlabel metal1 1644 1682 1756 1698 0 _1059_.gnd
rlabel metal1 1644 1442 1756 1458 0 _1059_.vdd
rlabel metal2 1653 1573 1667 1587 0 _1059_.A
rlabel metal2 1673 1553 1687 1567 0 _1059_.B
rlabel metal2 1693 1573 1707 1587 0 _1059_.C
rlabel metal2 1713 1553 1727 1567 0 _1059_.Y
rlabel metal1 2104 1682 2216 1698 0 _1005_.gnd
rlabel metal1 2104 1442 2216 1458 0 _1005_.vdd
rlabel metal2 2193 1593 2207 1607 0 _1005_.A
rlabel metal2 2173 1573 2187 1587 0 _1005_.B
rlabel metal2 2133 1573 2147 1587 0 _1005_.C
rlabel metal2 2153 1593 2167 1607 0 _1005_.Y
rlabel metal1 1944 1682 2016 1698 0 _1060_.gnd
rlabel metal1 1944 1442 2016 1458 0 _1060_.vdd
rlabel metal2 1953 1613 1967 1627 0 _1060_.A
rlabel metal2 1973 1573 1987 1587 0 _1060_.Y
rlabel metal1 2004 1682 2116 1698 0 _1004_.gnd
rlabel metal1 2004 1442 2116 1458 0 _1004_.vdd
rlabel metal2 2013 1573 2027 1587 0 _1004_.A
rlabel metal2 2033 1553 2047 1567 0 _1004_.B
rlabel metal2 2053 1573 2067 1587 0 _1004_.C
rlabel metal2 2073 1553 2087 1567 0 _1004_.Y
rlabel metal1 2264 1682 2516 1698 0 _1535_.gnd
rlabel metal1 2264 1442 2516 1458 0 _1535_.vdd
rlabel metal2 2413 1593 2427 1607 0 _1535_.D
rlabel metal2 2373 1593 2387 1607 0 _1535_.CLK
rlabel metal2 2293 1593 2307 1607 0 _1535_.Q
rlabel metal1 2204 1682 2276 1698 0 _953_.gnd
rlabel metal1 2204 1442 2276 1458 0 _953_.vdd
rlabel metal2 2213 1613 2227 1627 0 _953_.A
rlabel metal2 2233 1573 2247 1587 0 _953_.Y
rlabel metal1 2504 1682 2616 1698 0 _1369_.gnd
rlabel metal1 2504 1442 2616 1458 0 _1369_.vdd
rlabel metal2 2593 1593 2607 1607 0 _1369_.A
rlabel metal2 2573 1573 2587 1587 0 _1369_.B
rlabel metal2 2533 1573 2547 1587 0 _1369_.C
rlabel metal2 2553 1593 2567 1607 0 _1369_.Y
rlabel metal1 2604 1682 2716 1698 0 _1367_.gnd
rlabel metal1 2604 1442 2716 1458 0 _1367_.vdd
rlabel metal2 2693 1593 2707 1607 0 _1367_.A
rlabel metal2 2633 1593 2647 1607 0 _1367_.Y
rlabel metal2 2653 1553 2667 1567 0 _1367_.B
rlabel metal1 2784 1682 2896 1698 0 _1363_.gnd
rlabel metal1 2784 1442 2896 1458 0 _1363_.vdd
rlabel metal2 2793 1573 2807 1587 0 _1363_.A
rlabel metal2 2813 1613 2827 1627 0 _1363_.B
rlabel metal2 2833 1573 2847 1587 0 _1363_.C
rlabel metal2 2853 1593 2867 1607 0 _1363_.Y
rlabel metal1 2704 1682 2796 1698 0 _1368_.gnd
rlabel metal1 2704 1442 2796 1458 0 _1368_.vdd
rlabel metal2 2753 1593 2767 1607 0 _1368_.B
rlabel metal2 2713 1593 2727 1607 0 _1368_.A
rlabel metal2 2733 1613 2747 1627 0 _1368_.Y
rlabel metal1 2884 1682 2976 1698 0 _1354_.gnd
rlabel metal1 2884 1442 2976 1458 0 _1354_.vdd
rlabel metal2 2913 1593 2927 1607 0 _1354_.B
rlabel metal2 2953 1593 2967 1607 0 _1354_.A
rlabel metal2 2933 1613 2947 1627 0 _1354_.Y
rlabel metal1 3084 1682 3196 1698 0 _817_.gnd
rlabel metal1 3084 1442 3196 1458 0 _817_.vdd
rlabel metal2 3093 1593 3107 1607 0 _817_.A
rlabel metal2 3113 1573 3127 1587 0 _817_.B
rlabel metal2 3153 1573 3167 1587 0 _817_.C
rlabel metal2 3133 1593 3147 1607 0 _817_.Y
rlabel metal1 3184 1682 3276 1698 0 _816_.gnd
rlabel metal1 3184 1442 3276 1458 0 _816_.vdd
rlabel metal2 3193 1553 3207 1567 0 _816_.A
rlabel metal2 3233 1553 3247 1567 0 _816_.B
rlabel metal2 3213 1573 3227 1587 0 _816_.Y
rlabel metal1 2964 1682 3036 1698 0 _913_.gnd
rlabel metal1 2964 1442 3036 1458 0 _913_.vdd
rlabel metal2 3013 1613 3027 1627 0 _913_.A
rlabel metal2 2993 1573 3007 1587 0 _913_.Y
rlabel metal1 3024 1682 3096 1698 0 _815_.gnd
rlabel metal1 3024 1442 3096 1458 0 _815_.vdd
rlabel metal2 3073 1613 3087 1627 0 _815_.A
rlabel metal2 3053 1573 3067 1587 0 _815_.Y
rlabel metal1 3444 1682 3696 1698 0 _1565_.gnd
rlabel metal1 3444 1442 3696 1458 0 _1565_.vdd
rlabel metal2 3533 1593 3547 1607 0 _1565_.D
rlabel metal2 3573 1593 3587 1607 0 _1565_.CLK
rlabel metal2 3653 1593 3667 1607 0 _1565_.Q
rlabel metal1 3344 1682 3456 1698 0 _1370_.gnd
rlabel metal1 3344 1442 3456 1458 0 _1370_.vdd
rlabel metal2 3433 1593 3447 1607 0 _1370_.A
rlabel metal2 3413 1573 3427 1587 0 _1370_.B
rlabel metal2 3373 1573 3387 1587 0 _1370_.C
rlabel metal2 3393 1593 3407 1607 0 _1370_.Y
rlabel metal1 3264 1682 3356 1698 0 _810_.gnd
rlabel metal1 3264 1442 3356 1458 0 _810_.vdd
rlabel metal2 3333 1553 3347 1567 0 _810_.A
rlabel metal2 3293 1553 3307 1567 0 _810_.B
rlabel metal2 3313 1573 3327 1587 0 _810_.Y
rlabel metal1 3684 1682 3756 1698 0 _1362_.gnd
rlabel metal1 3684 1442 3756 1458 0 _1362_.vdd
rlabel metal2 3693 1613 3707 1627 0 _1362_.A
rlabel metal2 3713 1573 3727 1587 0 _1362_.Y
rlabel metal1 3804 1682 3916 1698 0 _1456_.gnd
rlabel metal1 3804 1442 3916 1458 0 _1456_.vdd
rlabel metal2 3893 1593 3907 1607 0 _1456_.A
rlabel metal2 3873 1573 3887 1587 0 _1456_.B
rlabel metal2 3833 1573 3847 1587 0 _1456_.C
rlabel metal2 3853 1593 3867 1607 0 _1456_.Y
rlabel metal1 3984 1682 4076 1698 0 _1449_.gnd
rlabel metal1 3984 1442 4076 1458 0 _1449_.vdd
rlabel metal2 4033 1593 4047 1607 0 _1449_.B
rlabel metal2 3993 1593 4007 1607 0 _1449_.A
rlabel metal2 4013 1613 4027 1627 0 _1449_.Y
rlabel metal1 3904 1682 3996 1698 0 _1448_.gnd
rlabel metal1 3904 1442 3996 1458 0 _1448_.vdd
rlabel metal2 3953 1593 3967 1607 0 _1448_.B
rlabel metal2 3913 1593 3927 1607 0 _1448_.A
rlabel metal2 3933 1613 3947 1627 0 _1448_.Y
rlabel metal1 3744 1682 3816 1698 0 _1455_.gnd
rlabel metal1 3744 1442 3816 1458 0 _1455_.vdd
rlabel metal2 3793 1613 3807 1627 0 _1455_.A
rlabel metal2 3773 1573 3787 1587 0 _1455_.Y
rlabel metal1 4124 1682 4236 1698 0 _1462_.gnd
rlabel metal1 4124 1442 4236 1458 0 _1462_.vdd
rlabel metal2 4133 1573 4147 1587 0 _1462_.A
rlabel metal2 4153 1613 4167 1627 0 _1462_.B
rlabel metal2 4173 1573 4187 1587 0 _1462_.C
rlabel metal2 4193 1593 4207 1607 0 _1462_.Y
rlabel metal1 4224 1682 4316 1698 0 _1466_.gnd
rlabel metal1 4224 1442 4316 1458 0 _1466_.vdd
rlabel metal2 4273 1593 4287 1607 0 _1466_.B
rlabel metal2 4233 1593 4247 1607 0 _1466_.A
rlabel metal2 4253 1613 4267 1627 0 _1466_.Y
rlabel metal1 4064 1682 4136 1698 0 _1451_.gnd
rlabel metal1 4064 1442 4136 1458 0 _1451_.vdd
rlabel metal2 4073 1613 4087 1627 0 _1451_.A
rlabel metal2 4093 1573 4107 1587 0 _1451_.Y
rlabel metal1 4304 1682 4416 1698 0 _1471_.gnd
rlabel metal1 4304 1442 4416 1458 0 _1471_.vdd
rlabel metal2 4313 1573 4327 1587 0 _1471_.A
rlabel metal2 4333 1613 4347 1627 0 _1471_.B
rlabel metal2 4353 1573 4367 1587 0 _1471_.C
rlabel metal2 4373 1593 4387 1607 0 _1471_.Y
rlabel metal1 4404 1682 4476 1698 0 _1470_.gnd
rlabel metal1 4404 1442 4476 1458 0 _1470_.vdd
rlabel metal2 4413 1613 4427 1627 0 _1470_.A
rlabel metal2 4433 1573 4447 1587 0 _1470_.Y
rlabel metal1 4464 1682 4536 1698 0 _1467_.gnd
rlabel metal1 4464 1442 4536 1458 0 _1467_.vdd
rlabel metal2 4473 1613 4487 1627 0 _1467_.A
rlabel metal2 4493 1573 4507 1587 0 _1467_.Y
rlabel metal1 4524 1682 4596 1698 0 _842_.gnd
rlabel metal1 4524 1442 4596 1458 0 _842_.vdd
rlabel metal2 4573 1613 4587 1627 0 _842_.A
rlabel metal2 4553 1573 4567 1587 0 _842_.Y
rlabel metal1 4584 1682 4696 1698 0 _1468_.gnd
rlabel metal1 4584 1442 4696 1458 0 _1468_.vdd
rlabel metal2 4593 1593 4607 1607 0 _1468_.A
rlabel metal2 4613 1573 4627 1587 0 _1468_.B
rlabel metal2 4653 1573 4667 1587 0 _1468_.C
rlabel metal2 4633 1593 4647 1607 0 _1468_.Y
rlabel metal1 4684 1682 4776 1698 0 _849_.gnd
rlabel metal1 4684 1442 4776 1458 0 _849_.vdd
rlabel metal2 4693 1553 4707 1567 0 _849_.A
rlabel metal2 4733 1553 4747 1567 0 _849_.B
rlabel metal2 4713 1573 4727 1587 0 _849_.Y
rlabel metal1 124 1682 236 1698 0 _1036_.gnd
rlabel metal1 124 1922 236 1938 0 _1036_.vdd
rlabel metal2 133 1773 147 1787 0 _1036_.A
rlabel metal2 153 1793 167 1807 0 _1036_.B
rlabel metal2 193 1793 207 1807 0 _1036_.C
rlabel metal2 173 1773 187 1787 0 _1036_.Y
rlabel metal1 224 1682 316 1698 0 _1030_.gnd
rlabel metal1 224 1922 316 1938 0 _1030_.vdd
rlabel metal2 233 1813 247 1827 0 _1030_.A
rlabel metal2 273 1813 287 1827 0 _1030_.B
rlabel metal2 253 1793 267 1807 0 _1030_.Y
rlabel metal1 4 1682 136 1698 0 _1089_.gnd
rlabel metal1 4 1922 136 1938 0 _1089_.vdd
rlabel metal2 113 1773 127 1787 0 _1089_.A
rlabel metal2 93 1793 107 1807 0 _1089_.B
rlabel metal2 33 1773 47 1787 0 _1089_.C
rlabel metal2 53 1793 67 1807 0 _1089_.D
rlabel metal2 73 1773 87 1787 0 _1089_.Y
rlabel metal1 304 1682 416 1698 0 _1031_.gnd
rlabel metal1 304 1922 416 1938 0 _1031_.vdd
rlabel metal2 393 1793 407 1807 0 _1031_.A
rlabel metal2 373 1813 387 1827 0 _1031_.B
rlabel metal2 353 1793 367 1807 0 _1031_.C
rlabel metal2 333 1813 347 1827 0 _1031_.Y
rlabel metal1 404 1682 536 1698 0 _1101_.gnd
rlabel metal1 404 1922 536 1938 0 _1101_.vdd
rlabel metal2 413 1773 427 1787 0 _1101_.A
rlabel metal2 433 1793 447 1807 0 _1101_.B
rlabel metal2 493 1773 507 1787 0 _1101_.C
rlabel metal2 473 1793 487 1807 0 _1101_.D
rlabel metal2 453 1773 467 1787 0 _1101_.Y
rlabel metal1 524 1682 636 1698 0 _1034_.gnd
rlabel metal1 524 1922 636 1938 0 _1034_.vdd
rlabel metal2 533 1773 547 1787 0 _1034_.A
rlabel metal2 593 1773 607 1787 0 _1034_.Y
rlabel metal2 573 1813 587 1827 0 _1034_.B
rlabel metal1 684 1682 776 1698 0 BUFX2_insert31.gnd
rlabel metal1 684 1922 776 1938 0 BUFX2_insert31.vdd
rlabel metal2 693 1773 707 1787 0 BUFX2_insert31.A
rlabel metal2 733 1773 747 1787 0 BUFX2_insert31.Y
rlabel metal1 764 1682 876 1698 0 _1120_.gnd
rlabel metal1 764 1922 876 1938 0 _1120_.vdd
rlabel metal2 853 1773 867 1787 0 _1120_.A
rlabel metal2 833 1793 847 1807 0 _1120_.B
rlabel metal2 793 1793 807 1807 0 _1120_.C
rlabel metal2 813 1773 827 1787 0 _1120_.Y
rlabel metal1 624 1682 696 1698 0 _860_.gnd
rlabel metal1 624 1922 696 1938 0 _860_.vdd
rlabel metal2 673 1793 687 1807 0 _860_.A
rlabel metal2 653 1773 667 1787 0 _860_.Y
rlabel metal1 864 1682 976 1698 0 _1116_.gnd
rlabel metal1 864 1922 976 1938 0 _1116_.vdd
rlabel metal2 873 1773 887 1787 0 _1116_.A
rlabel metal2 893 1793 907 1807 0 _1116_.B
rlabel metal2 933 1793 947 1807 0 _1116_.C
rlabel metal2 913 1773 927 1787 0 _1116_.Y
rlabel metal1 1064 1682 1136 1698 0 _1118_.gnd
rlabel metal1 1064 1922 1136 1938 0 _1118_.vdd
rlabel metal2 1073 1753 1087 1767 0 _1118_.A
rlabel metal2 1093 1793 1107 1807 0 _1118_.Y
rlabel metal1 964 1682 1076 1698 0 _1119_.gnd
rlabel metal1 964 1922 1076 1938 0 _1119_.vdd
rlabel metal2 973 1793 987 1807 0 _1119_.A
rlabel metal2 993 1813 1007 1827 0 _1119_.B
rlabel metal2 1013 1793 1027 1807 0 _1119_.C
rlabel metal2 1033 1813 1047 1827 0 _1119_.Y
rlabel metal1 1324 1682 1396 1698 0 _959_.gnd
rlabel metal1 1324 1922 1396 1938 0 _959_.vdd
rlabel metal2 1373 1753 1387 1767 0 _959_.A
rlabel metal2 1353 1793 1367 1807 0 _959_.Y
rlabel metal1 1224 1682 1336 1698 0 _1123_.gnd
rlabel metal1 1224 1922 1336 1938 0 _1123_.vdd
rlabel metal2 1233 1793 1247 1807 0 _1123_.A
rlabel metal2 1253 1813 1267 1827 0 _1123_.B
rlabel metal2 1273 1793 1287 1807 0 _1123_.C
rlabel metal2 1293 1813 1307 1827 0 _1123_.Y
rlabel metal1 1124 1682 1236 1698 0 _1121_.gnd
rlabel metal1 1124 1922 1236 1938 0 _1121_.vdd
rlabel metal2 1133 1793 1147 1807 0 _1121_.A
rlabel metal2 1153 1813 1167 1827 0 _1121_.B
rlabel metal2 1173 1793 1187 1807 0 _1121_.C
rlabel metal2 1193 1813 1207 1827 0 _1121_.Y
rlabel metal1 1604 1682 1676 1698 0 _1129_.gnd
rlabel metal1 1604 1922 1676 1938 0 _1129_.vdd
rlabel metal2 1613 1753 1627 1767 0 _1129_.A
rlabel metal2 1633 1793 1647 1807 0 _1129_.Y
rlabel metal1 1504 1682 1616 1698 0 _1130_.gnd
rlabel metal1 1504 1922 1616 1938 0 _1130_.vdd
rlabel metal2 1513 1793 1527 1807 0 _1130_.A
rlabel metal2 1533 1813 1547 1827 0 _1130_.B
rlabel metal2 1553 1793 1567 1807 0 _1130_.C
rlabel metal2 1573 1813 1587 1827 0 _1130_.Y
rlabel metal1 1384 1682 1516 1698 0 _1125_.gnd
rlabel metal1 1384 1922 1516 1938 0 _1125_.vdd
rlabel metal2 1493 1773 1507 1787 0 _1125_.A
rlabel metal2 1473 1793 1487 1807 0 _1125_.B
rlabel metal2 1413 1773 1427 1787 0 _1125_.C
rlabel metal2 1433 1793 1447 1807 0 _1125_.D
rlabel metal2 1453 1773 1467 1787 0 _1125_.Y
rlabel metal1 1724 1682 1836 1698 0 _1071_.gnd
rlabel metal1 1724 1922 1836 1938 0 _1071_.vdd
rlabel metal2 1813 1793 1827 1807 0 _1071_.A
rlabel metal2 1793 1813 1807 1827 0 _1071_.B
rlabel metal2 1773 1793 1787 1807 0 _1071_.C
rlabel metal2 1753 1813 1767 1827 0 _1071_.Y
rlabel metal1 1824 1682 1936 1698 0 _1065_.gnd
rlabel metal1 1824 1922 1936 1938 0 _1065_.vdd
rlabel metal2 1833 1773 1847 1787 0 _1065_.A
rlabel metal2 1893 1773 1907 1787 0 _1065_.Y
rlabel metal2 1873 1813 1887 1827 0 _1065_.B
rlabel metal1 1664 1682 1736 1698 0 _962_.gnd
rlabel metal1 1664 1922 1736 1938 0 _962_.vdd
rlabel metal2 1713 1793 1727 1807 0 _962_.A
rlabel metal2 1693 1773 1707 1787 0 _962_.Y
rlabel metal1 1924 1682 2176 1698 0 _1551_.gnd
rlabel metal1 1924 1922 2176 1938 0 _1551_.vdd
rlabel metal2 2013 1773 2027 1787 0 _1551_.D
rlabel metal2 2053 1773 2067 1787 0 _1551_.CLK
rlabel metal2 2133 1773 2147 1787 0 _1551_.Q
rlabel metal1 2304 1682 2416 1698 0 _820_.gnd
rlabel metal1 2304 1922 2416 1938 0 _820_.vdd
rlabel metal2 2313 1773 2327 1787 0 _820_.A
rlabel metal2 2333 1793 2347 1807 0 _820_.B
rlabel metal2 2373 1793 2387 1807 0 _820_.C
rlabel metal2 2353 1773 2367 1787 0 _820_.Y
rlabel metal1 2404 1682 2496 1698 0 _1366_.gnd
rlabel metal1 2404 1922 2496 1938 0 _1366_.vdd
rlabel metal2 2453 1773 2467 1787 0 _1366_.B
rlabel metal2 2413 1773 2427 1787 0 _1366_.A
rlabel metal2 2433 1753 2447 1767 0 _1366_.Y
rlabel metal1 2164 1682 2256 1698 0 _1364_.gnd
rlabel metal1 2164 1922 2256 1938 0 _1364_.vdd
rlabel metal2 2193 1773 2207 1787 0 _1364_.B
rlabel metal2 2233 1773 2247 1787 0 _1364_.A
rlabel metal2 2213 1753 2227 1767 0 _1364_.Y
rlabel metal1 2244 1682 2316 1698 0 _818_.gnd
rlabel metal1 2244 1922 2316 1938 0 _818_.vdd
rlabel metal2 2253 1753 2267 1767 0 _818_.A
rlabel metal2 2273 1793 2287 1807 0 _818_.Y
rlabel metal1 2564 1682 2676 1698 0 _1373_.gnd
rlabel metal1 2564 1922 2676 1938 0 _1373_.vdd
rlabel metal2 2573 1773 2587 1787 0 _1373_.A
rlabel metal2 2593 1793 2607 1807 0 _1373_.B
rlabel metal2 2633 1793 2647 1807 0 _1373_.C
rlabel metal2 2613 1773 2627 1787 0 _1373_.Y
rlabel metal1 2664 1682 2756 1698 0 _1372_.gnd
rlabel metal1 2664 1922 2756 1938 0 _1372_.vdd
rlabel metal2 2733 1813 2747 1827 0 _1372_.A
rlabel metal2 2693 1813 2707 1827 0 _1372_.B
rlabel metal2 2713 1793 2727 1807 0 _1372_.Y
rlabel metal1 2484 1682 2576 1698 0 _1365_.gnd
rlabel metal1 2484 1922 2576 1938 0 _1365_.vdd
rlabel metal2 2533 1773 2547 1787 0 _1365_.B
rlabel metal2 2493 1773 2507 1787 0 _1365_.A
rlabel metal2 2513 1753 2527 1767 0 _1365_.Y
rlabel metal1 2824 1682 2936 1698 0 _1357_.gnd
rlabel metal1 2824 1922 2936 1938 0 _1357_.vdd
rlabel metal2 2833 1773 2847 1787 0 _1357_.A
rlabel metal2 2853 1793 2867 1807 0 _1357_.B
rlabel metal2 2893 1793 2907 1807 0 _1357_.C
rlabel metal2 2873 1773 2887 1787 0 _1357_.Y
rlabel metal1 2744 1682 2836 1698 0 _1358_.gnd
rlabel metal1 2744 1922 2836 1938 0 _1358_.vdd
rlabel metal2 2773 1773 2787 1787 0 _1358_.B
rlabel metal2 2813 1773 2827 1787 0 _1358_.A
rlabel metal2 2793 1753 2807 1767 0 _1358_.Y
rlabel metal1 2924 1682 2996 1698 0 _1356_.gnd
rlabel metal1 2924 1922 2996 1938 0 _1356_.vdd
rlabel metal2 2933 1753 2947 1767 0 _1356_.A
rlabel metal2 2953 1793 2967 1807 0 _1356_.Y
rlabel metal1 3064 1682 3316 1698 0 _1534_.gnd
rlabel metal1 3064 1922 3316 1938 0 _1534_.vdd
rlabel metal2 3213 1773 3227 1787 0 _1534_.D
rlabel metal2 3173 1773 3187 1787 0 _1534_.CLK
rlabel metal2 3093 1773 3107 1787 0 _1534_.Q
rlabel metal1 2984 1682 3076 1698 0 _1353_.gnd
rlabel metal1 2984 1922 3076 1938 0 _1353_.vdd
rlabel metal2 3013 1773 3027 1787 0 _1353_.B
rlabel metal2 3053 1773 3067 1787 0 _1353_.A
rlabel metal2 3033 1753 3047 1767 0 _1353_.Y
rlabel metal1 3304 1682 3416 1698 0 _1351_.gnd
rlabel metal1 3304 1922 3416 1938 0 _1351_.vdd
rlabel metal2 3313 1773 3327 1787 0 _1351_.A
rlabel metal2 3333 1793 3347 1807 0 _1351_.B
rlabel metal2 3373 1793 3387 1807 0 _1351_.C
rlabel metal2 3353 1773 3367 1787 0 _1351_.Y
rlabel metal1 3404 1682 3496 1698 0 _1350_.gnd
rlabel metal1 3404 1922 3496 1938 0 _1350_.vdd
rlabel metal2 3413 1813 3427 1827 0 _1350_.A
rlabel metal2 3453 1813 3467 1827 0 _1350_.B
rlabel metal2 3433 1793 3447 1807 0 _1350_.Y
rlabel metal1 3724 1682 3816 1698 0 BUFX2_insert16.gnd
rlabel metal1 3724 1922 3816 1938 0 BUFX2_insert16.vdd
rlabel metal2 3733 1773 3747 1787 0 BUFX2_insert16.A
rlabel metal2 3773 1773 3787 1787 0 BUFX2_insert16.Y
rlabel metal1 3484 1682 3736 1698 0 _1563_.gnd
rlabel metal1 3484 1922 3736 1938 0 _1563_.vdd
rlabel metal2 3633 1773 3647 1787 0 _1563_.D
rlabel metal2 3593 1773 3607 1787 0 _1563_.CLK
rlabel metal2 3513 1773 3527 1787 0 _1563_.Q
rlabel metal1 3884 1682 3996 1698 0 _1453_.gnd
rlabel metal1 3884 1922 3996 1938 0 _1453_.vdd
rlabel metal2 3973 1773 3987 1787 0 _1453_.A
rlabel metal2 3953 1793 3967 1807 0 _1453_.B
rlabel metal2 3913 1793 3927 1807 0 _1453_.C
rlabel metal2 3933 1773 3947 1787 0 _1453_.Y
rlabel metal1 3984 1682 4096 1698 0 _1452_.gnd
rlabel metal1 3984 1922 4096 1938 0 _1452_.vdd
rlabel metal2 4073 1773 4087 1787 0 _1452_.A
rlabel metal2 4053 1793 4067 1807 0 _1452_.B
rlabel metal2 4013 1793 4027 1807 0 _1452_.C
rlabel metal2 4033 1773 4047 1787 0 _1452_.Y
rlabel metal1 3804 1682 3896 1698 0 _1438_.gnd
rlabel metal1 3804 1922 3896 1938 0 _1438_.vdd
rlabel metal2 3873 1813 3887 1827 0 _1438_.A
rlabel metal2 3833 1813 3847 1827 0 _1438_.B
rlabel metal2 3853 1793 3867 1807 0 _1438_.Y
rlabel metal1 4244 1682 4356 1698 0 _1465_.gnd
rlabel metal1 4244 1922 4356 1938 0 _1465_.vdd
rlabel metal2 4253 1793 4267 1807 0 _1465_.A
rlabel metal2 4273 1753 4287 1767 0 _1465_.B
rlabel metal2 4293 1793 4307 1807 0 _1465_.C
rlabel metal2 4313 1773 4327 1787 0 _1465_.Y
rlabel metal1 4184 1682 4256 1698 0 _1460_.gnd
rlabel metal1 4184 1922 4256 1938 0 _1460_.vdd
rlabel metal2 4233 1753 4247 1767 0 _1460_.A
rlabel metal2 4213 1793 4227 1807 0 _1460_.Y
rlabel metal1 4084 1682 4196 1698 0 _1461_.gnd
rlabel metal1 4084 1922 4196 1938 0 _1461_.vdd
rlabel metal2 4093 1753 4107 1767 0 _1461_.A
rlabel metal2 4113 1773 4127 1787 0 _1461_.B
rlabel metal2 4153 1793 4167 1807 0 _1461_.Y
rlabel metal1 4424 1682 4676 1698 0 _1574_.gnd
rlabel metal1 4424 1922 4676 1938 0 _1574_.vdd
rlabel metal2 4573 1773 4587 1787 0 _1574_.D
rlabel metal2 4533 1773 4547 1787 0 _1574_.CLK
rlabel metal2 4453 1773 4467 1787 0 _1574_.Q
rlabel metal1 4344 1682 4436 1698 0 _1459_.gnd
rlabel metal1 4344 1922 4436 1938 0 _1459_.vdd
rlabel metal2 4373 1773 4387 1787 0 _1459_.B
rlabel metal2 4413 1773 4427 1787 0 _1459_.A
rlabel metal2 4393 1753 4407 1767 0 _1459_.Y
rlabel nsubstratencontact 4756 1928 4756 1928 0 FILL71250x25350.vdd
rlabel metal1 4744 1682 4776 1698 0 FILL71250x25350.gnd
rlabel metal1 4664 1682 4756 1698 0 _846_.gnd
rlabel metal1 4664 1922 4756 1938 0 _846_.vdd
rlabel metal2 4733 1813 4747 1827 0 _846_.A
rlabel metal2 4693 1813 4707 1827 0 _846_.B
rlabel metal2 4713 1793 4727 1807 0 _846_.Y
rlabel metal1 4 2162 96 2178 0 BUFX2_insert33.gnd
rlabel metal1 4 1922 96 1938 0 BUFX2_insert33.vdd
rlabel metal2 73 2073 87 2087 0 BUFX2_insert33.A
rlabel metal2 33 2073 47 2087 0 BUFX2_insert33.Y
rlabel metal1 84 2162 196 2178 0 _1029_.gnd
rlabel metal1 84 1922 196 1938 0 _1029_.vdd
rlabel metal2 173 2073 187 2087 0 _1029_.A
rlabel metal2 153 2053 167 2067 0 _1029_.B
rlabel metal2 113 2053 127 2067 0 _1029_.C
rlabel metal2 133 2073 147 2087 0 _1029_.Y
rlabel metal1 184 2162 296 2178 0 _1106_.gnd
rlabel metal1 184 1922 296 1938 0 _1106_.vdd
rlabel metal2 273 2053 287 2067 0 _1106_.A
rlabel metal2 253 2033 267 2047 0 _1106_.B
rlabel metal2 233 2053 247 2067 0 _1106_.C
rlabel metal2 213 2033 227 2047 0 _1106_.Y
rlabel metal1 284 2162 396 2178 0 _1115_.gnd
rlabel metal1 284 1922 396 1938 0 _1115_.vdd
rlabel metal2 293 2053 307 2067 0 _1115_.A
rlabel metal2 313 2093 327 2107 0 _1115_.B
rlabel metal2 333 2053 347 2067 0 _1115_.C
rlabel metal2 353 2073 367 2087 0 _1115_.Y
rlabel metal1 384 2162 496 2178 0 _1114_.gnd
rlabel metal1 384 1922 496 1938 0 _1114_.vdd
rlabel metal2 393 2053 407 2067 0 _1114_.A
rlabel metal2 413 2093 427 2107 0 _1114_.B
rlabel metal2 433 2053 447 2067 0 _1114_.C
rlabel metal2 453 2073 467 2087 0 _1114_.Y
rlabel metal1 484 2162 596 2178 0 _1110_.gnd
rlabel metal1 484 1922 596 1938 0 _1110_.vdd
rlabel metal2 493 2053 507 2067 0 _1110_.A
rlabel metal2 513 2033 527 2047 0 _1110_.B
rlabel metal2 533 2053 547 2067 0 _1110_.C
rlabel metal2 553 2033 567 2047 0 _1110_.Y
rlabel metal1 784 2162 896 2178 0 _1141_.gnd
rlabel metal1 784 1922 896 1938 0 _1141_.vdd
rlabel metal2 873 2073 887 2087 0 _1141_.A
rlabel metal2 853 2053 867 2067 0 _1141_.B
rlabel metal2 813 2053 827 2067 0 _1141_.C
rlabel metal2 833 2073 847 2087 0 _1141_.Y
rlabel metal1 684 2162 796 2178 0 _1140_.gnd
rlabel metal1 684 1922 796 1938 0 _1140_.vdd
rlabel metal2 693 2053 707 2067 0 _1140_.A
rlabel metal2 713 2093 727 2107 0 _1140_.B
rlabel metal2 733 2053 747 2067 0 _1140_.C
rlabel metal2 753 2073 767 2087 0 _1140_.Y
rlabel metal1 584 2162 696 2178 0 _1111_.gnd
rlabel metal1 584 1922 696 1938 0 _1111_.vdd
rlabel metal2 593 2053 607 2067 0 _1111_.A
rlabel metal2 613 2033 627 2047 0 _1111_.B
rlabel metal2 633 2053 647 2067 0 _1111_.C
rlabel metal2 653 2033 667 2047 0 _1111_.Y
rlabel metal1 884 2162 996 2178 0 _1124_.gnd
rlabel metal1 884 1922 996 1938 0 _1124_.vdd
rlabel metal2 893 2053 907 2067 0 _1124_.A
rlabel metal2 913 2033 927 2047 0 _1124_.B
rlabel metal2 933 2053 947 2067 0 _1124_.C
rlabel metal2 953 2033 967 2047 0 _1124_.Y
rlabel metal1 984 2162 1096 2178 0 _1117_.gnd
rlabel metal1 984 1922 1096 1938 0 _1117_.vdd
rlabel metal2 993 2053 1007 2067 0 _1117_.A
rlabel metal2 1013 2033 1027 2047 0 _1117_.B
rlabel metal2 1033 2053 1047 2067 0 _1117_.C
rlabel metal2 1053 2033 1067 2047 0 _1117_.Y
rlabel metal1 1184 2162 1296 2178 0 _1122_.gnd
rlabel metal1 1184 1922 1296 1938 0 _1122_.vdd
rlabel metal2 1193 2053 1207 2067 0 _1122_.A
rlabel metal2 1213 2093 1227 2107 0 _1122_.B
rlabel metal2 1233 2053 1247 2067 0 _1122_.C
rlabel metal2 1253 2073 1267 2087 0 _1122_.Y
rlabel metal1 1284 2162 1376 2178 0 _1126_.gnd
rlabel metal1 1284 1922 1376 1938 0 _1126_.vdd
rlabel metal2 1333 2073 1347 2087 0 _1126_.B
rlabel metal2 1293 2073 1307 2087 0 _1126_.A
rlabel metal2 1313 2093 1327 2107 0 _1126_.Y
rlabel metal1 1084 2162 1196 2178 0 _1131_.gnd
rlabel metal1 1084 1922 1196 1938 0 _1131_.vdd
rlabel metal2 1093 2053 1107 2067 0 _1131_.A
rlabel metal2 1113 2033 1127 2047 0 _1131_.B
rlabel metal2 1133 2053 1147 2067 0 _1131_.C
rlabel metal2 1153 2033 1167 2047 0 _1131_.Y
rlabel metal1 1604 2162 1716 2178 0 _1139_.gnd
rlabel metal1 1604 1922 1716 1938 0 _1139_.vdd
rlabel metal2 1693 2073 1707 2087 0 _1139_.A
rlabel metal2 1673 2053 1687 2067 0 _1139_.B
rlabel metal2 1633 2053 1647 2067 0 _1139_.C
rlabel metal2 1653 2073 1667 2087 0 _1139_.Y
rlabel metal1 1444 2162 1536 2178 0 _1138_.gnd
rlabel metal1 1444 1922 1536 1938 0 _1138_.vdd
rlabel metal2 1513 2033 1527 2047 0 _1138_.A
rlabel metal2 1473 2033 1487 2047 0 _1138_.B
rlabel metal2 1493 2053 1507 2067 0 _1138_.Y
rlabel metal1 1364 2162 1456 2178 0 _1137_.gnd
rlabel metal1 1364 1922 1456 1938 0 _1137_.vdd
rlabel metal2 1433 2033 1447 2047 0 _1137_.A
rlabel metal2 1393 2033 1407 2047 0 _1137_.B
rlabel metal2 1413 2053 1427 2067 0 _1137_.Y
rlabel metal1 1524 2162 1616 2178 0 _1132_.gnd
rlabel metal1 1524 1922 1616 1938 0 _1132_.vdd
rlabel metal2 1533 2033 1547 2047 0 _1132_.A
rlabel metal2 1573 2033 1587 2047 0 _1132_.B
rlabel metal2 1553 2053 1567 2067 0 _1132_.Y
rlabel metal1 1704 2162 1816 2178 0 _1127_.gnd
rlabel metal1 1704 1922 1816 1938 0 _1127_.vdd
rlabel metal2 1713 2053 1727 2067 0 _1127_.A
rlabel metal2 1733 2093 1747 2107 0 _1127_.B
rlabel metal2 1753 2053 1767 2067 0 _1127_.C
rlabel metal2 1773 2073 1787 2087 0 _1127_.Y
rlabel metal1 1804 2162 1896 2178 0 _1133_.gnd
rlabel metal1 1804 1922 1896 1938 0 _1133_.vdd
rlabel metal2 1853 2073 1867 2087 0 _1133_.B
rlabel metal2 1813 2073 1827 2087 0 _1133_.A
rlabel metal2 1833 2093 1847 2107 0 _1133_.Y
rlabel metal1 2084 2162 2196 2178 0 _1135_.gnd
rlabel metal1 2084 1922 2196 1938 0 _1135_.vdd
rlabel metal2 2173 2073 2187 2087 0 _1135_.A
rlabel metal2 2153 2053 2167 2067 0 _1135_.B
rlabel metal2 2113 2053 2127 2067 0 _1135_.C
rlabel metal2 2133 2073 2147 2087 0 _1135_.Y
rlabel metal1 1984 2162 2096 2178 0 _1134_.gnd
rlabel metal1 1984 1922 2096 1938 0 _1134_.vdd
rlabel metal2 1993 2073 2007 2087 0 _1134_.A
rlabel metal2 2013 2053 2027 2067 0 _1134_.B
rlabel metal2 2053 2053 2067 2067 0 _1134_.C
rlabel metal2 2033 2073 2047 2087 0 _1134_.Y
rlabel metal1 1884 2162 1996 2178 0 _1128_.gnd
rlabel metal1 1884 1922 1996 1938 0 _1128_.vdd
rlabel metal2 1973 2073 1987 2087 0 _1128_.A
rlabel metal2 1953 2053 1967 2067 0 _1128_.B
rlabel metal2 1913 2053 1927 2067 0 _1128_.C
rlabel metal2 1933 2073 1947 2087 0 _1128_.Y
rlabel metal1 2184 2162 2396 2178 0 CLKBUF1_insert11.gnd
rlabel metal1 2184 1922 2396 1938 0 CLKBUF1_insert11.vdd
rlabel metal2 2353 2053 2367 2067 0 CLKBUF1_insert11.A
rlabel metal2 2213 2053 2227 2067 0 CLKBUF1_insert11.Y
rlabel metal1 2384 2162 2476 2178 0 _819_.gnd
rlabel metal1 2384 1922 2476 1938 0 _819_.vdd
rlabel metal2 2393 2033 2407 2047 0 _819_.A
rlabel metal2 2433 2033 2447 2047 0 _819_.B
rlabel metal2 2413 2053 2427 2067 0 _819_.Y
rlabel metal1 2664 2162 2756 2178 0 _1359_.gnd
rlabel metal1 2664 1922 2756 1938 0 _1359_.vdd
rlabel metal2 2733 2033 2747 2047 0 _1359_.A
rlabel metal2 2693 2033 2707 2047 0 _1359_.B
rlabel metal2 2713 2053 2727 2067 0 _1359_.Y
rlabel metal1 2564 2162 2676 2178 0 _1313_.gnd
rlabel metal1 2564 1922 2676 1938 0 _1313_.vdd
rlabel metal2 2573 2093 2587 2107 0 _1313_.A
rlabel metal2 2593 2073 2607 2087 0 _1313_.B
rlabel metal2 2633 2053 2647 2067 0 _1313_.Y
rlabel metal1 2464 2162 2576 2178 0 _1374_.gnd
rlabel metal1 2464 1922 2576 1938 0 _1374_.vdd
rlabel metal2 2553 2073 2567 2087 0 _1374_.A
rlabel metal2 2493 2073 2507 2087 0 _1374_.Y
rlabel metal2 2513 2033 2527 2047 0 _1374_.B
rlabel metal1 2824 2162 3076 2178 0 _1589_.gnd
rlabel metal1 2824 1922 3076 1938 0 _1589_.vdd
rlabel metal2 2913 2073 2927 2087 0 _1589_.D
rlabel metal2 2953 2073 2967 2087 0 _1589_.CLK
rlabel metal2 3033 2073 3047 2087 0 _1589_.Q
rlabel metal1 2744 2162 2836 2178 0 _1360_.gnd
rlabel metal1 2744 1922 2836 1938 0 _1360_.vdd
rlabel metal2 2753 2033 2767 2047 0 _1360_.A
rlabel metal2 2793 2033 2807 2047 0 _1360_.B
rlabel metal2 2773 2053 2787 2067 0 _1360_.Y
rlabel metal1 3064 2162 3176 2178 0 _1513_.gnd
rlabel metal1 3064 1922 3176 1938 0 _1513_.vdd
rlabel metal2 3153 2053 3167 2067 0 _1513_.A
rlabel metal2 3133 2093 3147 2107 0 _1513_.B
rlabel metal2 3113 2053 3127 2067 0 _1513_.C
rlabel metal2 3093 2073 3107 2087 0 _1513_.Y
rlabel metal1 3164 2162 3256 2178 0 _1512_.gnd
rlabel metal1 3164 1922 3256 1938 0 _1512_.vdd
rlabel metal2 3213 2073 3227 2087 0 _1512_.B
rlabel metal2 3173 2073 3187 2087 0 _1512_.A
rlabel metal2 3193 2093 3207 2107 0 _1512_.Y
rlabel metal1 3364 2162 3616 2178 0 _1559_.gnd
rlabel metal1 3364 1922 3616 1938 0 _1559_.vdd
rlabel metal2 3453 2073 3467 2087 0 _1559_.D
rlabel metal2 3493 2073 3507 2087 0 _1559_.CLK
rlabel metal2 3573 2073 3587 2087 0 _1559_.Q
rlabel metal1 3244 2162 3376 2178 0 _1317_.gnd
rlabel metal1 3244 1922 3376 1938 0 _1317_.vdd
rlabel metal2 3353 2073 3367 2087 0 _1317_.A
rlabel metal2 3333 2053 3347 2067 0 _1317_.B
rlabel metal2 3273 2073 3287 2087 0 _1317_.C
rlabel metal2 3293 2053 3307 2067 0 _1317_.D
rlabel metal2 3313 2073 3327 2087 0 _1317_.Y
rlabel metal1 3704 2162 3956 2178 0 _1564_.gnd
rlabel metal1 3704 1922 3956 1938 0 _1564_.vdd
rlabel metal2 3793 2073 3807 2087 0 _1564_.D
rlabel metal2 3833 2073 3847 2087 0 _1564_.CLK
rlabel metal2 3913 2073 3927 2087 0 _1564_.Q
rlabel metal1 3604 2162 3716 2178 0 _1361_.gnd
rlabel metal1 3604 1922 3716 1938 0 _1361_.vdd
rlabel metal2 3613 2073 3627 2087 0 _1361_.A
rlabel metal2 3633 2053 3647 2067 0 _1361_.B
rlabel metal2 3673 2053 3687 2067 0 _1361_.C
rlabel metal2 3653 2073 3667 2087 0 _1361_.Y
rlabel metal1 3944 2162 4196 2178 0 _1572_.gnd
rlabel metal1 3944 1922 4196 1938 0 _1572_.vdd
rlabel metal2 4093 2073 4107 2087 0 _1572_.D
rlabel metal2 4053 2073 4067 2087 0 _1572_.CLK
rlabel metal2 3973 2073 3987 2087 0 _1572_.Q
rlabel metal1 4184 2162 4316 2178 0 _1463_.gnd
rlabel metal1 4184 1922 4316 1938 0 _1463_.vdd
rlabel metal2 4293 2073 4307 2087 0 _1463_.A
rlabel metal2 4273 2053 4287 2067 0 _1463_.B
rlabel metal2 4213 2073 4227 2087 0 _1463_.C
rlabel metal2 4233 2053 4247 2067 0 _1463_.D
rlabel metal2 4253 2073 4267 2087 0 _1463_.Y
rlabel metal1 4524 2162 4776 2178 0 _1543_.gnd
rlabel metal1 4524 1922 4776 1938 0 _1543_.vdd
rlabel metal2 4673 2073 4687 2087 0 _1543_.D
rlabel metal2 4633 2073 4647 2087 0 _1543_.CLK
rlabel metal2 4553 2073 4567 2087 0 _1543_.Q
rlabel metal1 4364 2162 4456 2178 0 _1458_.gnd
rlabel metal1 4364 1922 4456 1938 0 _1458_.vdd
rlabel metal2 4393 2073 4407 2087 0 _1458_.B
rlabel metal2 4433 2073 4447 2087 0 _1458_.A
rlabel metal2 4413 2093 4427 2107 0 _1458_.Y
rlabel metal1 4444 2162 4536 2178 0 _1457_.gnd
rlabel metal1 4444 1922 4536 1938 0 _1457_.vdd
rlabel metal2 4473 2073 4487 2087 0 _1457_.B
rlabel metal2 4513 2073 4527 2087 0 _1457_.A
rlabel metal2 4493 2093 4507 2107 0 _1457_.Y
rlabel metal1 4304 2162 4376 2178 0 _1312_.gnd
rlabel metal1 4304 1922 4376 1938 0 _1312_.vdd
rlabel metal2 4313 2093 4327 2107 0 _1312_.A
rlabel metal2 4333 2053 4347 2067 0 _1312_.Y
rlabel metal1 104 2162 216 2178 0 _1109_.gnd
rlabel metal1 104 2402 216 2418 0 _1109_.vdd
rlabel metal2 193 2253 207 2267 0 _1109_.A
rlabel metal2 173 2273 187 2287 0 _1109_.B
rlabel metal2 133 2273 147 2287 0 _1109_.C
rlabel metal2 153 2253 167 2267 0 _1109_.Y
rlabel metal1 204 2162 316 2178 0 _1105_.gnd
rlabel metal1 204 2402 316 2418 0 _1105_.vdd
rlabel metal2 213 2253 227 2267 0 _1105_.A
rlabel metal2 233 2273 247 2287 0 _1105_.B
rlabel metal2 273 2273 287 2287 0 _1105_.C
rlabel metal2 253 2253 267 2267 0 _1105_.Y
rlabel metal1 4 2162 116 2178 0 _1100_.gnd
rlabel metal1 4 2402 116 2418 0 _1100_.vdd
rlabel metal2 93 2273 107 2287 0 _1100_.A
rlabel metal2 73 2293 87 2307 0 _1100_.B
rlabel metal2 53 2273 67 2287 0 _1100_.C
rlabel metal2 33 2293 47 2307 0 _1100_.Y
rlabel metal1 504 2162 616 2178 0 _1177_.gnd
rlabel metal1 504 2402 616 2418 0 _1177_.vdd
rlabel metal2 513 2253 527 2267 0 _1177_.A
rlabel metal2 533 2273 547 2287 0 _1177_.B
rlabel metal2 573 2273 587 2287 0 _1177_.C
rlabel metal2 553 2253 567 2267 0 _1177_.Y
rlabel metal1 404 2162 516 2178 0 _1176_.gnd
rlabel metal1 404 2402 516 2418 0 _1176_.vdd
rlabel metal2 413 2273 427 2287 0 _1176_.A
rlabel metal2 433 2233 447 2247 0 _1176_.B
rlabel metal2 453 2273 467 2287 0 _1176_.C
rlabel metal2 473 2253 487 2267 0 _1176_.Y
rlabel metal1 304 2162 416 2178 0 _1108_.gnd
rlabel metal1 304 2402 416 2418 0 _1108_.vdd
rlabel metal2 313 2273 327 2287 0 _1108_.A
rlabel metal2 333 2293 347 2307 0 _1108_.B
rlabel metal2 353 2273 367 2287 0 _1108_.C
rlabel metal2 373 2293 387 2307 0 _1108_.Y
rlabel metal1 604 2162 716 2178 0 _1145_.gnd
rlabel metal1 604 2402 716 2418 0 _1145_.vdd
rlabel metal2 693 2273 707 2287 0 _1145_.A
rlabel metal2 673 2233 687 2247 0 _1145_.B
rlabel metal2 653 2273 667 2287 0 _1145_.C
rlabel metal2 633 2253 647 2267 0 _1145_.Y
rlabel metal1 704 2162 776 2178 0 _1144_.gnd
rlabel metal1 704 2402 776 2418 0 _1144_.vdd
rlabel metal2 713 2233 727 2247 0 _1144_.A
rlabel metal2 733 2273 747 2287 0 _1144_.Y
rlabel metal1 764 2162 876 2178 0 _1107_.gnd
rlabel metal1 764 2402 876 2418 0 _1107_.vdd
rlabel metal2 853 2253 867 2267 0 _1107_.A
rlabel metal2 793 2253 807 2267 0 _1107_.Y
rlabel metal2 813 2293 827 2307 0 _1107_.B
rlabel metal1 1044 2162 1156 2178 0 _1079_.gnd
rlabel metal1 1044 2402 1156 2418 0 _1079_.vdd
rlabel metal2 1133 2253 1147 2267 0 _1079_.A
rlabel metal2 1113 2273 1127 2287 0 _1079_.B
rlabel metal2 1073 2273 1087 2287 0 _1079_.C
rlabel metal2 1093 2253 1107 2267 0 _1079_.Y
rlabel metal1 864 2162 956 2178 0 _1088_.gnd
rlabel metal1 864 2402 956 2418 0 _1088_.vdd
rlabel metal2 873 2293 887 2307 0 _1088_.A
rlabel metal2 913 2293 927 2307 0 _1088_.B
rlabel metal2 893 2273 907 2287 0 _1088_.Y
rlabel metal1 944 2162 1056 2178 0 _1078_.gnd
rlabel metal1 944 2402 1056 2418 0 _1078_.vdd
rlabel metal2 953 2253 967 2267 0 _1078_.A
rlabel metal2 1013 2253 1027 2267 0 _1078_.Y
rlabel metal2 993 2293 1007 2307 0 _1078_.B
rlabel metal1 1244 2162 1496 2178 0 _1594_.gnd
rlabel metal1 1244 2402 1496 2418 0 _1594_.vdd
rlabel metal2 1333 2253 1347 2267 0 _1594_.D
rlabel metal2 1373 2253 1387 2267 0 _1594_.CLK
rlabel metal2 1453 2253 1467 2267 0 _1594_.Q
rlabel metal1 1144 2162 1256 2178 0 _1523_.gnd
rlabel metal1 1144 2402 1256 2418 0 _1523_.vdd
rlabel metal2 1233 2253 1247 2267 0 _1523_.A
rlabel metal2 1213 2273 1227 2287 0 _1523_.B
rlabel metal2 1173 2273 1187 2287 0 _1523_.C
rlabel metal2 1193 2253 1207 2267 0 _1523_.Y
rlabel metal1 1584 2162 1836 2178 0 _1592_.gnd
rlabel metal1 1584 2402 1836 2418 0 _1592_.vdd
rlabel metal2 1673 2253 1687 2267 0 _1592_.D
rlabel metal2 1713 2253 1727 2267 0 _1592_.CLK
rlabel metal2 1793 2253 1807 2267 0 _1592_.Q
rlabel metal1 1484 2162 1596 2178 0 _1519_.gnd
rlabel metal1 1484 2402 1596 2418 0 _1519_.vdd
rlabel metal2 1573 2253 1587 2267 0 _1519_.A
rlabel metal2 1553 2273 1567 2287 0 _1519_.B
rlabel metal2 1513 2273 1527 2287 0 _1519_.C
rlabel metal2 1533 2253 1547 2267 0 _1519_.Y
rlabel metal1 1824 2162 1896 2178 0 _1003_.gnd
rlabel metal1 1824 2402 1896 2418 0 _1003_.vdd
rlabel metal2 1873 2233 1887 2247 0 _1003_.A
rlabel metal2 1853 2273 1867 2287 0 _1003_.Y
rlabel metal1 2044 2162 2296 2178 0 _1553_.gnd
rlabel metal1 2044 2402 2296 2418 0 _1553_.vdd
rlabel metal2 2133 2253 2147 2267 0 _1553_.D
rlabel metal2 2173 2253 2187 2267 0 _1553_.CLK
rlabel metal2 2253 2253 2267 2267 0 _1553_.Q
rlabel metal1 1944 2162 2056 2178 0 _1068_.gnd
rlabel metal1 1944 2402 2056 2418 0 _1068_.vdd
rlabel metal2 1953 2253 1967 2267 0 _1068_.A
rlabel metal2 1973 2273 1987 2287 0 _1068_.B
rlabel metal2 2013 2273 2027 2287 0 _1068_.C
rlabel metal2 1993 2253 2007 2267 0 _1068_.Y
rlabel metal1 1884 2162 1956 2178 0 _1067_.gnd
rlabel metal1 1884 2402 1956 2418 0 _1067_.vdd
rlabel metal2 1933 2233 1947 2247 0 _1067_.A
rlabel metal2 1913 2273 1927 2287 0 _1067_.Y
rlabel metal1 2284 2162 2396 2178 0 _1397_.gnd
rlabel metal1 2284 2402 2396 2418 0 _1397_.vdd
rlabel metal2 2373 2273 2387 2287 0 _1397_.A
rlabel metal2 2353 2233 2367 2247 0 _1397_.B
rlabel metal2 2333 2273 2347 2287 0 _1397_.C
rlabel metal2 2313 2253 2327 2267 0 _1397_.Y
rlabel metal1 2384 2162 2496 2178 0 _1375_.gnd
rlabel metal1 2384 2402 2496 2418 0 _1375_.vdd
rlabel metal2 2473 2273 2487 2287 0 _1375_.A
rlabel metal2 2453 2233 2467 2247 0 _1375_.B
rlabel metal2 2433 2273 2447 2287 0 _1375_.C
rlabel metal2 2413 2253 2427 2267 0 _1375_.Y
rlabel metal1 2484 2162 2596 2178 0 _1398_.gnd
rlabel metal1 2484 2402 2596 2418 0 _1398_.vdd
rlabel metal2 2493 2273 2507 2287 0 _1398_.A
rlabel metal2 2513 2293 2527 2307 0 _1398_.B
rlabel metal2 2533 2273 2547 2287 0 _1398_.C
rlabel metal2 2553 2293 2567 2307 0 _1398_.Y
rlabel metal1 2584 2162 2696 2178 0 _1399_.gnd
rlabel metal1 2584 2402 2696 2418 0 _1399_.vdd
rlabel metal2 2593 2253 2607 2267 0 _1399_.A
rlabel metal2 2653 2253 2667 2267 0 _1399_.Y
rlabel metal2 2633 2293 2647 2307 0 _1399_.B
rlabel metal1 2684 2162 2936 2178 0 _1585_.gnd
rlabel metal1 2684 2402 2936 2418 0 _1585_.vdd
rlabel metal2 2833 2253 2847 2267 0 _1585_.D
rlabel metal2 2793 2253 2807 2267 0 _1585_.CLK
rlabel metal2 2713 2253 2727 2267 0 _1585_.Q
rlabel metal1 2924 2162 3036 2178 0 _1504_.gnd
rlabel metal1 2924 2402 3036 2418 0 _1504_.vdd
rlabel metal2 3013 2253 3027 2267 0 _1504_.A
rlabel metal2 2993 2273 3007 2287 0 _1504_.B
rlabel metal2 2953 2273 2967 2287 0 _1504_.C
rlabel metal2 2973 2253 2987 2267 0 _1504_.Y
rlabel metal1 3024 2162 3136 2178 0 _1505_.gnd
rlabel metal1 3024 2402 3136 2418 0 _1505_.vdd
rlabel metal2 3113 2253 3127 2267 0 _1505_.A
rlabel metal2 3093 2273 3107 2287 0 _1505_.B
rlabel metal2 3053 2273 3067 2287 0 _1505_.C
rlabel metal2 3073 2253 3087 2267 0 _1505_.Y
rlabel metal1 3124 2162 3236 2178 0 _1502_.gnd
rlabel metal1 3124 2402 3236 2418 0 _1502_.vdd
rlabel metal2 3133 2253 3147 2267 0 _1502_.A
rlabel metal2 3153 2273 3167 2287 0 _1502_.B
rlabel metal2 3193 2273 3207 2287 0 _1502_.C
rlabel metal2 3173 2253 3187 2267 0 _1502_.Y
rlabel metal1 3224 2162 3476 2178 0 _1584_.gnd
rlabel metal1 3224 2402 3476 2418 0 _1584_.vdd
rlabel metal2 3373 2253 3387 2267 0 _1584_.D
rlabel metal2 3333 2253 3347 2267 0 _1584_.CLK
rlabel metal2 3253 2253 3267 2267 0 _1584_.Q
rlabel metal1 3464 2162 3576 2178 0 _1503_.gnd
rlabel metal1 3464 2402 3576 2418 0 _1503_.vdd
rlabel metal2 3553 2253 3567 2267 0 _1503_.A
rlabel metal2 3533 2273 3547 2287 0 _1503_.B
rlabel metal2 3493 2273 3507 2287 0 _1503_.C
rlabel metal2 3513 2253 3527 2267 0 _1503_.Y
rlabel metal1 3564 2162 3656 2178 0 _1450_.gnd
rlabel metal1 3564 2402 3656 2418 0 _1450_.vdd
rlabel metal2 3593 2253 3607 2267 0 _1450_.B
rlabel metal2 3633 2253 3647 2267 0 _1450_.A
rlabel metal2 3613 2233 3627 2247 0 _1450_.Y
rlabel metal1 3644 2162 3756 2178 0 _1445_.gnd
rlabel metal1 3644 2402 3756 2418 0 _1445_.vdd
rlabel metal2 3653 2233 3667 2247 0 _1445_.A
rlabel metal2 3673 2253 3687 2267 0 _1445_.B
rlabel metal2 3713 2273 3727 2287 0 _1445_.Y
rlabel metal1 3744 2162 3836 2178 0 _1352_.gnd
rlabel metal1 3744 2402 3836 2418 0 _1352_.vdd
rlabel metal2 3813 2293 3827 2307 0 _1352_.A
rlabel metal2 3773 2293 3787 2307 0 _1352_.B
rlabel metal2 3793 2273 3807 2287 0 _1352_.Y
rlabel metal1 3824 2162 3956 2178 0 _772_.gnd
rlabel metal1 3824 2402 3956 2418 0 _772_.vdd
rlabel metal2 3933 2253 3947 2267 0 _772_.A
rlabel metal2 3913 2273 3927 2287 0 _772_.B
rlabel metal2 3853 2253 3867 2267 0 _772_.C
rlabel metal2 3873 2273 3887 2287 0 _772_.D
rlabel metal2 3893 2253 3907 2267 0 _772_.Y
rlabel metal1 3944 2162 4076 2178 0 _766_.gnd
rlabel metal1 3944 2402 4076 2418 0 _766_.vdd
rlabel metal2 4053 2253 4067 2267 0 _766_.A
rlabel metal2 4033 2273 4047 2287 0 _766_.B
rlabel metal2 3973 2253 3987 2267 0 _766_.C
rlabel metal2 3993 2273 4007 2287 0 _766_.D
rlabel metal2 4013 2253 4027 2267 0 _766_.Y
rlabel metal1 4064 2162 4316 2178 0 _1573_.gnd
rlabel metal1 4064 2402 4316 2418 0 _1573_.vdd
rlabel metal2 4153 2253 4167 2267 0 _1573_.D
rlabel metal2 4193 2253 4207 2267 0 _1573_.CLK
rlabel metal2 4273 2253 4287 2267 0 _1573_.Q
rlabel metal1 4304 2162 4556 2178 0 _1576_.gnd
rlabel metal1 4304 2402 4556 2418 0 _1576_.vdd
rlabel metal2 4453 2253 4467 2267 0 _1576_.D
rlabel metal2 4413 2253 4427 2267 0 _1576_.CLK
rlabel metal2 4333 2253 4347 2267 0 _1576_.Q
rlabel nsubstratencontact 4756 2408 4756 2408 0 FILL71250x32550.vdd
rlabel metal1 4744 2162 4776 2178 0 FILL71250x32550.gnd
rlabel nsubstratencontact 4736 2408 4736 2408 0 FILL70950x32550.vdd
rlabel metal1 4724 2162 4756 2178 0 FILL70950x32550.gnd
rlabel metal1 4544 2162 4656 2178 0 _1482_.gnd
rlabel metal1 4544 2402 4656 2418 0 _1482_.vdd
rlabel metal2 4553 2253 4567 2267 0 _1482_.A
rlabel metal2 4573 2273 4587 2287 0 _1482_.B
rlabel metal2 4613 2273 4627 2287 0 _1482_.C
rlabel metal2 4593 2253 4607 2267 0 _1482_.Y
rlabel metal1 4644 2162 4736 2178 0 _1481_.gnd
rlabel metal1 4644 2402 4736 2418 0 _1481_.vdd
rlabel metal2 4653 2293 4667 2307 0 _1481_.A
rlabel metal2 4693 2293 4707 2307 0 _1481_.B
rlabel metal2 4673 2273 4687 2287 0 _1481_.Y
rlabel metal1 104 2642 216 2658 0 _1103_.gnd
rlabel metal1 104 2402 216 2418 0 _1103_.vdd
rlabel metal2 113 2533 127 2547 0 _1103_.A
rlabel metal2 133 2573 147 2587 0 _1103_.B
rlabel metal2 153 2533 167 2547 0 _1103_.C
rlabel metal2 173 2553 187 2567 0 _1103_.Y
rlabel metal1 204 2642 276 2658 0 _1095_.gnd
rlabel metal1 204 2402 276 2418 0 _1095_.vdd
rlabel metal2 253 2573 267 2587 0 _1095_.A
rlabel metal2 233 2533 247 2547 0 _1095_.Y
rlabel metal1 4 2642 116 2658 0 _1099_.gnd
rlabel metal1 4 2402 116 2418 0 _1099_.vdd
rlabel metal2 13 2533 27 2547 0 _1099_.A
rlabel metal2 33 2513 47 2527 0 _1099_.B
rlabel metal2 53 2533 67 2547 0 _1099_.C
rlabel metal2 73 2513 87 2527 0 _1099_.Y
rlabel metal1 264 2642 376 2658 0 _1028_.gnd
rlabel metal1 264 2402 376 2418 0 _1028_.vdd
rlabel metal2 353 2553 367 2567 0 _1028_.A
rlabel metal2 293 2553 307 2567 0 _1028_.Y
rlabel metal2 313 2513 327 2527 0 _1028_.B
rlabel metal1 364 2642 476 2658 0 _1104_.gnd
rlabel metal1 364 2402 476 2418 0 _1104_.vdd
rlabel metal2 453 2533 467 2547 0 _1104_.A
rlabel metal2 433 2573 447 2587 0 _1104_.B
rlabel metal2 413 2533 427 2547 0 _1104_.C
rlabel metal2 393 2553 407 2567 0 _1104_.Y
rlabel metal1 464 2642 576 2658 0 _1094_.gnd
rlabel metal1 464 2402 576 2418 0 _1094_.vdd
rlabel metal2 553 2533 567 2547 0 _1094_.A
rlabel metal2 533 2513 547 2527 0 _1094_.B
rlabel metal2 513 2533 527 2547 0 _1094_.C
rlabel metal2 493 2513 507 2527 0 _1094_.Y
rlabel metal1 564 2642 676 2658 0 _1093_.gnd
rlabel metal1 564 2402 676 2418 0 _1093_.vdd
rlabel metal2 653 2553 667 2567 0 _1093_.A
rlabel metal2 633 2533 647 2547 0 _1093_.B
rlabel metal2 593 2533 607 2547 0 _1093_.C
rlabel metal2 613 2553 627 2567 0 _1093_.Y
rlabel metal1 724 2642 816 2658 0 _1142_.gnd
rlabel metal1 724 2402 816 2418 0 _1142_.vdd
rlabel metal2 793 2513 807 2527 0 _1142_.A
rlabel metal2 753 2513 767 2527 0 _1142_.B
rlabel metal2 773 2533 787 2547 0 _1142_.Y
rlabel metal1 664 2642 736 2658 0 _899_.gnd
rlabel metal1 664 2402 736 2418 0 _899_.vdd
rlabel metal2 713 2533 727 2547 0 _899_.A
rlabel metal2 693 2553 707 2567 0 _899_.Y
rlabel metal1 904 2642 1016 2658 0 _1086_.gnd
rlabel metal1 904 2402 1016 2418 0 _1086_.vdd
rlabel metal2 993 2553 1007 2567 0 _1086_.A
rlabel metal2 973 2533 987 2547 0 _1086_.B
rlabel metal2 933 2533 947 2547 0 _1086_.C
rlabel metal2 953 2553 967 2567 0 _1086_.Y
rlabel metal1 1004 2642 1096 2658 0 _1084_.gnd
rlabel metal1 1004 2402 1096 2418 0 _1084_.vdd
rlabel metal2 1013 2513 1027 2527 0 _1084_.A
rlabel metal2 1053 2513 1067 2527 0 _1084_.B
rlabel metal2 1033 2533 1047 2547 0 _1084_.Y
rlabel metal1 804 2642 916 2658 0 _1087_.gnd
rlabel metal1 804 2402 916 2418 0 _1087_.vdd
rlabel metal2 893 2533 907 2547 0 _1087_.A
rlabel metal2 873 2513 887 2527 0 _1087_.B
rlabel metal2 853 2533 867 2547 0 _1087_.C
rlabel metal2 833 2513 847 2527 0 _1087_.Y
rlabel metal1 1244 2642 1356 2658 0 _1521_.gnd
rlabel metal1 1244 2402 1356 2418 0 _1521_.vdd
rlabel metal2 1333 2553 1347 2567 0 _1521_.A
rlabel metal2 1313 2533 1327 2547 0 _1521_.B
rlabel metal2 1273 2533 1287 2547 0 _1521_.C
rlabel metal2 1293 2553 1307 2567 0 _1521_.Y
rlabel metal1 1184 2642 1256 2658 0 _1083_.gnd
rlabel metal1 1184 2402 1256 2418 0 _1083_.vdd
rlabel metal2 1233 2573 1247 2587 0 _1083_.A
rlabel metal2 1213 2533 1227 2547 0 _1083_.Y
rlabel metal1 1084 2642 1196 2658 0 _1082_.gnd
rlabel metal1 1084 2402 1196 2418 0 _1082_.vdd
rlabel metal2 1173 2533 1187 2547 0 _1082_.A
rlabel metal2 1153 2513 1167 2527 0 _1082_.B
rlabel metal2 1133 2533 1147 2547 0 _1082_.C
rlabel metal2 1113 2513 1127 2527 0 _1082_.Y
rlabel metal1 1564 2642 1816 2658 0 _1593_.gnd
rlabel metal1 1564 2402 1816 2418 0 _1593_.vdd
rlabel metal2 1653 2553 1667 2567 0 _1593_.D
rlabel metal2 1693 2553 1707 2567 0 _1593_.CLK
rlabel metal2 1773 2553 1787 2567 0 _1593_.Q
rlabel metal1 1484 2642 1576 2658 0 _1518_.gnd
rlabel metal1 1484 2402 1576 2418 0 _1518_.vdd
rlabel metal2 1553 2513 1567 2527 0 _1518_.A
rlabel metal2 1513 2513 1527 2527 0 _1518_.B
rlabel metal2 1533 2533 1547 2547 0 _1518_.Y
rlabel metal1 1344 2642 1436 2658 0 _1077_.gnd
rlabel metal1 1344 2402 1436 2418 0 _1077_.vdd
rlabel metal2 1353 2513 1367 2527 0 _1077_.A
rlabel metal2 1393 2513 1407 2527 0 _1077_.B
rlabel metal2 1373 2533 1387 2547 0 _1077_.Y
rlabel metal1 1424 2642 1496 2658 0 _786_.gnd
rlabel metal1 1424 2402 1496 2418 0 _786_.vdd
rlabel metal2 1433 2533 1447 2547 0 _786_.A
rlabel metal2 1453 2553 1467 2567 0 _786_.Y
rlabel metal1 1804 2642 1896 2658 0 _784_.gnd
rlabel metal1 1804 2402 1896 2418 0 _784_.vdd
rlabel metal2 1813 2513 1827 2527 0 _784_.A
rlabel metal2 1853 2513 1867 2527 0 _784_.B
rlabel metal2 1833 2533 1847 2547 0 _784_.Y
rlabel metal1 1884 2642 1976 2658 0 _787_.gnd
rlabel metal1 1884 2402 1976 2418 0 _787_.vdd
rlabel metal2 1893 2513 1907 2527 0 _787_.A
rlabel metal2 1933 2513 1947 2527 0 _787_.B
rlabel metal2 1913 2533 1927 2547 0 _787_.Y
rlabel metal1 2064 2642 2156 2658 0 _1066_.gnd
rlabel metal1 2064 2402 2156 2418 0 _1066_.vdd
rlabel metal2 2113 2553 2127 2567 0 _1066_.B
rlabel metal2 2073 2553 2087 2567 0 _1066_.A
rlabel metal2 2093 2573 2107 2587 0 _1066_.Y
rlabel metal1 1964 2642 2076 2658 0 _1269_.gnd
rlabel metal1 1964 2402 2076 2418 0 _1269_.vdd
rlabel metal2 1973 2533 1987 2547 0 _1269_.A
rlabel metal2 1993 2513 2007 2527 0 _1269_.B
rlabel metal2 2013 2533 2027 2547 0 _1269_.C
rlabel metal2 2033 2513 2047 2527 0 _1269_.Y
rlabel metal1 2344 2642 2456 2658 0 _1395_.gnd
rlabel metal1 2344 2402 2456 2418 0 _1395_.vdd
rlabel metal2 2433 2553 2447 2567 0 _1395_.A
rlabel metal2 2413 2533 2427 2547 0 _1395_.B
rlabel metal2 2373 2533 2387 2547 0 _1395_.C
rlabel metal2 2393 2553 2407 2567 0 _1395_.Y
rlabel metal1 2204 2642 2296 2658 0 _1386_.gnd
rlabel metal1 2204 2402 2296 2418 0 _1386_.vdd
rlabel metal2 2233 2553 2247 2567 0 _1386_.B
rlabel metal2 2273 2553 2287 2567 0 _1386_.A
rlabel metal2 2253 2573 2267 2587 0 _1386_.Y
rlabel metal1 2284 2642 2356 2658 0 _1394_.gnd
rlabel metal1 2284 2402 2356 2418 0 _1394_.vdd
rlabel metal2 2333 2573 2347 2587 0 _1394_.A
rlabel metal2 2313 2533 2327 2547 0 _1394_.Y
rlabel metal1 2144 2642 2216 2658 0 _1070_.gnd
rlabel metal1 2144 2402 2216 2418 0 _1070_.vdd
rlabel metal2 2193 2573 2207 2587 0 _1070_.A
rlabel metal2 2173 2533 2187 2547 0 _1070_.Y
rlabel metal1 2624 2642 2736 2658 0 _1384_.gnd
rlabel metal1 2624 2402 2736 2418 0 _1384_.vdd
rlabel metal2 2633 2553 2647 2567 0 _1384_.A
rlabel metal2 2653 2533 2667 2547 0 _1384_.B
rlabel metal2 2693 2533 2707 2547 0 _1384_.C
rlabel metal2 2673 2553 2687 2567 0 _1384_.Y
rlabel metal1 2444 2642 2536 2658 0 _1387_.gnd
rlabel metal1 2444 2402 2536 2418 0 _1387_.vdd
rlabel metal2 2493 2553 2507 2567 0 _1387_.B
rlabel metal2 2453 2553 2467 2567 0 _1387_.A
rlabel metal2 2473 2573 2487 2587 0 _1387_.Y
rlabel metal1 2524 2642 2636 2658 0 _1396_.gnd
rlabel metal1 2524 2402 2636 2418 0 _1396_.vdd
rlabel metal2 2533 2553 2547 2567 0 _1396_.A
rlabel metal2 2593 2553 2607 2567 0 _1396_.Y
rlabel metal2 2573 2513 2587 2527 0 _1396_.B
rlabel metal1 2904 2642 2996 2658 0 _1390_.gnd
rlabel metal1 2904 2402 2996 2418 0 _1390_.vdd
rlabel metal2 2913 2513 2927 2527 0 _1390_.A
rlabel metal2 2953 2513 2967 2527 0 _1390_.B
rlabel metal2 2933 2533 2947 2547 0 _1390_.Y
rlabel metal1 2724 2642 2816 2658 0 _1389_.gnd
rlabel metal1 2724 2402 2816 2418 0 _1389_.vdd
rlabel metal2 2793 2513 2807 2527 0 _1389_.A
rlabel metal2 2753 2513 2767 2527 0 _1389_.B
rlabel metal2 2773 2533 2787 2547 0 _1389_.Y
rlabel metal1 2804 2642 2916 2658 0 _1388_.gnd
rlabel metal1 2804 2402 2916 2418 0 _1388_.vdd
rlabel metal2 2813 2573 2827 2587 0 _1388_.A
rlabel metal2 2833 2553 2847 2567 0 _1388_.B
rlabel metal2 2873 2533 2887 2547 0 _1388_.Y
rlabel metal1 2984 2642 3076 2658 0 BUFX2_insert27.gnd
rlabel metal1 2984 2402 3076 2418 0 BUFX2_insert27.vdd
rlabel metal2 2993 2553 3007 2567 0 BUFX2_insert27.A
rlabel metal2 3033 2553 3047 2567 0 BUFX2_insert27.Y
rlabel metal1 3164 2642 3256 2658 0 BUFX2_insert19.gnd
rlabel metal1 3164 2402 3256 2418 0 BUFX2_insert19.vdd
rlabel metal2 3233 2553 3247 2567 0 BUFX2_insert19.A
rlabel metal2 3193 2553 3207 2567 0 BUFX2_insert19.Y
rlabel metal1 3064 2642 3176 2658 0 _1392_.gnd
rlabel metal1 3064 2402 3176 2418 0 _1392_.vdd
rlabel metal2 3073 2553 3087 2567 0 _1392_.A
rlabel metal2 3093 2533 3107 2547 0 _1392_.B
rlabel metal2 3133 2533 3147 2547 0 _1392_.C
rlabel metal2 3113 2553 3127 2567 0 _1392_.Y
rlabel metal1 3444 2642 3536 2658 0 BUFX2_insert28.gnd
rlabel metal1 3444 2402 3536 2418 0 BUFX2_insert28.vdd
rlabel metal2 3453 2553 3467 2567 0 BUFX2_insert28.A
rlabel metal2 3493 2553 3507 2567 0 BUFX2_insert28.Y
rlabel metal1 3244 2642 3336 2658 0 _1391_.gnd
rlabel metal1 3244 2402 3336 2418 0 _1391_.vdd
rlabel metal2 3313 2513 3327 2527 0 _1391_.A
rlabel metal2 3273 2513 3287 2527 0 _1391_.B
rlabel metal2 3293 2533 3307 2547 0 _1391_.Y
rlabel metal1 3324 2642 3456 2658 0 _781_.gnd
rlabel metal1 3324 2402 3456 2418 0 _781_.vdd
rlabel metal2 3333 2553 3347 2567 0 _781_.A
rlabel metal2 3353 2533 3367 2547 0 _781_.B
rlabel metal2 3413 2553 3427 2567 0 _781_.C
rlabel metal2 3393 2533 3407 2547 0 _781_.D
rlabel metal2 3373 2553 3387 2567 0 _781_.Y
rlabel metal1 3524 2642 3616 2658 0 BUFX2_insert17.gnd
rlabel metal1 3524 2402 3616 2418 0 BUFX2_insert17.vdd
rlabel metal2 3593 2553 3607 2567 0 BUFX2_insert17.A
rlabel metal2 3553 2553 3567 2567 0 BUFX2_insert17.Y
rlabel metal1 3604 2642 3856 2658 0 _1588_.gnd
rlabel metal1 3604 2402 3856 2418 0 _1588_.vdd
rlabel metal2 3693 2553 3707 2567 0 _1588_.D
rlabel metal2 3733 2553 3747 2567 0 _1588_.CLK
rlabel metal2 3813 2553 3827 2567 0 _1588_.Q
rlabel metal1 3844 2642 3956 2658 0 _1511_.gnd
rlabel metal1 3844 2402 3956 2418 0 _1511_.vdd
rlabel metal2 3933 2533 3947 2547 0 _1511_.A
rlabel metal2 3913 2573 3927 2587 0 _1511_.B
rlabel metal2 3893 2533 3907 2547 0 _1511_.C
rlabel metal2 3873 2553 3887 2567 0 _1511_.Y
rlabel metal1 3944 2642 4036 2658 0 _1510_.gnd
rlabel metal1 3944 2402 4036 2418 0 _1510_.vdd
rlabel metal2 3993 2553 4007 2567 0 _1510_.B
rlabel metal2 3953 2553 3967 2567 0 _1510_.A
rlabel metal2 3973 2573 3987 2587 0 _1510_.Y
rlabel metal1 4024 2642 4236 2658 0 CLKBUF1_insert14.gnd
rlabel metal1 4024 2402 4236 2418 0 CLKBUF1_insert14.vdd
rlabel metal2 4053 2533 4067 2547 0 CLKBUF1_insert14.A
rlabel metal2 4193 2533 4207 2547 0 CLKBUF1_insert14.Y
rlabel metal1 4224 2642 4476 2658 0 _1579_.gnd
rlabel metal1 4224 2402 4476 2418 0 _1579_.vdd
rlabel metal2 4313 2553 4327 2567 0 _1579_.D
rlabel metal2 4353 2553 4367 2567 0 _1579_.CLK
rlabel metal2 4433 2553 4447 2567 0 _1579_.Q
rlabel metal1 4464 2642 4576 2658 0 _1491_.gnd
rlabel metal1 4464 2402 4576 2418 0 _1491_.vdd
rlabel metal2 4473 2553 4487 2567 0 _1491_.A
rlabel metal2 4493 2533 4507 2547 0 _1491_.B
rlabel metal2 4533 2533 4547 2547 0 _1491_.C
rlabel metal2 4513 2553 4527 2567 0 _1491_.Y
rlabel nsubstratencontact 4764 2412 4764 2412 0 FILL71250x36150.vdd
rlabel metal1 4744 2642 4776 2658 0 FILL71250x36150.gnd
rlabel nsubstratencontact 4744 2412 4744 2412 0 FILL70950x36150.vdd
rlabel metal1 4724 2642 4756 2658 0 FILL70950x36150.gnd
rlabel metal1 4564 2642 4656 2658 0 _1490_.gnd
rlabel metal1 4564 2402 4656 2418 0 _1490_.vdd
rlabel metal2 4573 2513 4587 2527 0 _1490_.A
rlabel metal2 4613 2513 4627 2527 0 _1490_.B
rlabel metal2 4593 2533 4607 2547 0 _1490_.Y
rlabel metal1 4644 2642 4736 2658 0 _843_.gnd
rlabel metal1 4644 2402 4736 2418 0 _843_.vdd
rlabel metal2 4653 2513 4667 2527 0 _843_.A
rlabel metal2 4693 2513 4707 2527 0 _843_.B
rlabel metal2 4673 2533 4687 2547 0 _843_.Y
rlabel metal1 64 2642 176 2658 0 _1165_.gnd
rlabel metal1 64 2882 176 2898 0 _1165_.vdd
rlabel metal2 153 2733 167 2747 0 _1165_.A
rlabel metal2 133 2753 147 2767 0 _1165_.B
rlabel metal2 93 2753 107 2767 0 _1165_.C
rlabel metal2 113 2733 127 2747 0 _1165_.Y
rlabel metal1 4 2642 76 2658 0 _1098_.gnd
rlabel metal1 4 2882 76 2898 0 _1098_.vdd
rlabel metal2 53 2713 67 2727 0 _1098_.A
rlabel metal2 33 2753 47 2767 0 _1098_.Y
rlabel metal1 164 2642 296 2658 0 _1097_.gnd
rlabel metal1 164 2882 296 2898 0 _1097_.vdd
rlabel metal2 173 2733 187 2747 0 _1097_.A
rlabel metal2 193 2753 207 2767 0 _1097_.B
rlabel metal2 253 2733 267 2747 0 _1097_.C
rlabel metal2 233 2753 247 2767 0 _1097_.D
rlabel metal2 213 2733 227 2747 0 _1097_.Y
rlabel metal1 464 2642 576 2658 0 _1092_.gnd
rlabel metal1 464 2882 576 2898 0 _1092_.vdd
rlabel metal2 553 2733 567 2747 0 _1092_.A
rlabel metal2 533 2753 547 2767 0 _1092_.B
rlabel metal2 493 2753 507 2767 0 _1092_.C
rlabel metal2 513 2733 527 2747 0 _1092_.Y
rlabel metal1 284 2642 376 2658 0 _1096_.gnd
rlabel metal1 284 2882 376 2898 0 _1096_.vdd
rlabel metal2 293 2773 307 2787 0 _1096_.A
rlabel metal2 333 2773 347 2787 0 _1096_.B
rlabel metal2 313 2753 327 2767 0 _1096_.Y
rlabel metal1 364 2642 476 2658 0 _1091_.gnd
rlabel metal1 364 2882 476 2898 0 _1091_.vdd
rlabel metal2 373 2733 387 2747 0 _1091_.A
rlabel metal2 433 2733 447 2747 0 _1091_.Y
rlabel metal2 413 2773 427 2787 0 _1091_.B
rlabel metal1 564 2642 656 2658 0 _1090_.gnd
rlabel metal1 564 2882 656 2898 0 _1090_.vdd
rlabel metal2 573 2773 587 2787 0 _1090_.A
rlabel metal2 613 2773 627 2787 0 _1090_.B
rlabel metal2 593 2753 607 2767 0 _1090_.Y
rlabel metal1 764 2642 856 2658 0 _1085_.gnd
rlabel metal1 764 2882 856 2898 0 _1085_.vdd
rlabel metal2 773 2773 787 2787 0 _1085_.A
rlabel metal2 813 2773 827 2787 0 _1085_.B
rlabel metal2 793 2753 807 2767 0 _1085_.Y
rlabel metal1 644 2642 716 2658 0 _792_.gnd
rlabel metal1 644 2882 716 2898 0 _792_.vdd
rlabel metal2 693 2753 707 2767 0 _792_.A
rlabel metal2 673 2733 687 2747 0 _792_.Y
rlabel metal1 704 2642 776 2658 0 _783_.gnd
rlabel metal1 704 2882 776 2898 0 _783_.vdd
rlabel metal2 753 2753 767 2767 0 _783_.A
rlabel metal2 733 2733 747 2747 0 _783_.Y
rlabel metal1 944 2642 1056 2658 0 _1081_.gnd
rlabel metal1 944 2882 1056 2898 0 _1081_.vdd
rlabel metal2 1033 2733 1047 2747 0 _1081_.A
rlabel metal2 1013 2753 1027 2767 0 _1081_.B
rlabel metal2 973 2753 987 2767 0 _1081_.C
rlabel metal2 993 2733 1007 2747 0 _1081_.Y
rlabel metal1 1044 2642 1136 2658 0 _795_.gnd
rlabel metal1 1044 2882 1136 2898 0 _795_.vdd
rlabel metal2 1053 2773 1067 2787 0 _795_.A
rlabel metal2 1093 2773 1107 2787 0 _795_.B
rlabel metal2 1073 2753 1087 2767 0 _795_.Y
rlabel metal1 844 2642 956 2658 0 _1080_.gnd
rlabel metal1 844 2882 956 2898 0 _1080_.vdd
rlabel metal2 853 2733 867 2747 0 _1080_.A
rlabel metal2 913 2733 927 2747 0 _1080_.Y
rlabel metal2 893 2773 907 2787 0 _1080_.B
rlabel metal1 1224 2642 1476 2658 0 _1526_.gnd
rlabel metal1 1224 2882 1476 2898 0 _1526_.vdd
rlabel metal2 1373 2733 1387 2747 0 _1526_.D
rlabel metal2 1333 2733 1347 2747 0 _1526_.CLK
rlabel metal2 1253 2733 1267 2747 0 _1526_.Q
rlabel metal1 1124 2642 1236 2658 0 _796_.gnd
rlabel metal1 1124 2882 1236 2898 0 _796_.vdd
rlabel metal2 1213 2733 1227 2747 0 _796_.A
rlabel metal2 1193 2753 1207 2767 0 _796_.B
rlabel metal2 1153 2753 1167 2767 0 _796_.C
rlabel metal2 1173 2733 1187 2747 0 _796_.Y
rlabel metal1 1464 2642 1556 2658 0 BUFX2_insert29.gnd
rlabel metal1 1464 2882 1556 2898 0 BUFX2_insert29.vdd
rlabel metal2 1533 2733 1547 2747 0 BUFX2_insert29.A
rlabel metal2 1493 2733 1507 2747 0 BUFX2_insert29.Y
rlabel metal1 1544 2642 1796 2658 0 _1552_.gnd
rlabel metal1 1544 2882 1796 2898 0 _1552_.vdd
rlabel metal2 1633 2733 1647 2747 0 _1552_.D
rlabel metal2 1673 2733 1687 2747 0 _1552_.CLK
rlabel metal2 1753 2733 1767 2747 0 _1552_.Q
rlabel metal1 1784 2642 1896 2658 0 _788_.gnd
rlabel metal1 1784 2882 1896 2898 0 _788_.vdd
rlabel metal2 1793 2733 1807 2747 0 _788_.A
rlabel metal2 1813 2753 1827 2767 0 _788_.B
rlabel metal2 1853 2753 1867 2767 0 _788_.C
rlabel metal2 1833 2733 1847 2747 0 _788_.Y
rlabel metal1 2064 2642 2156 2658 0 _1376_.gnd
rlabel metal1 2064 2882 2156 2898 0 _1376_.vdd
rlabel metal2 2093 2733 2107 2747 0 _1376_.B
rlabel metal2 2133 2733 2147 2747 0 _1376_.A
rlabel metal2 2113 2713 2127 2727 0 _1376_.Y
rlabel metal1 1884 2642 1956 2658 0 _1006_.gnd
rlabel metal1 1884 2882 1956 2898 0 _1006_.vdd
rlabel metal2 1893 2713 1907 2727 0 _1006_.A
rlabel metal2 1913 2753 1927 2767 0 _1006_.Y
rlabel metal1 1944 2642 2076 2658 0 _1069_.gnd
rlabel metal1 1944 2882 2076 2898 0 _1069_.vdd
rlabel metal2 1953 2733 1967 2747 0 _1069_.A
rlabel metal2 1973 2753 1987 2767 0 _1069_.B
rlabel metal2 2033 2733 2047 2747 0 _1069_.C
rlabel metal2 1993 2733 2007 2747 0 _1069_.Y
rlabel metal2 2013 2753 2027 2767 0 _1069_.D
rlabel metal1 2364 2642 2456 2658 0 _1385_.gnd
rlabel metal1 2364 2882 2456 2898 0 _1385_.vdd
rlabel metal2 2393 2733 2407 2747 0 _1385_.B
rlabel metal2 2433 2733 2447 2747 0 _1385_.A
rlabel metal2 2413 2713 2427 2727 0 _1385_.Y
rlabel metal1 2224 2642 2316 2658 0 _1378_.gnd
rlabel metal1 2224 2882 2316 2898 0 _1378_.vdd
rlabel metal2 2253 2733 2267 2747 0 _1378_.B
rlabel metal2 2293 2733 2307 2747 0 _1378_.A
rlabel metal2 2273 2713 2287 2727 0 _1378_.Y
rlabel metal1 2144 2642 2236 2658 0 _1377_.gnd
rlabel metal1 2144 2882 2236 2898 0 _1377_.vdd
rlabel metal2 2173 2733 2187 2747 0 _1377_.B
rlabel metal2 2213 2733 2227 2747 0 _1377_.A
rlabel metal2 2193 2713 2207 2727 0 _1377_.Y
rlabel metal1 2304 2642 2376 2658 0 _1383_.gnd
rlabel metal1 2304 2882 2376 2898 0 _1383_.vdd
rlabel metal2 2313 2713 2327 2727 0 _1383_.A
rlabel metal2 2333 2753 2347 2767 0 _1383_.Y
rlabel metal1 2604 2642 2716 2658 0 _1381_.gnd
rlabel metal1 2604 2882 2716 2898 0 _1381_.vdd
rlabel metal2 2613 2733 2627 2747 0 _1381_.A
rlabel metal2 2633 2753 2647 2767 0 _1381_.B
rlabel metal2 2673 2753 2687 2767 0 _1381_.C
rlabel metal2 2653 2733 2667 2747 0 _1381_.Y
rlabel metal1 2444 2642 2516 2658 0 _1379_.gnd
rlabel metal1 2444 2882 2516 2898 0 _1379_.vdd
rlabel metal2 2453 2713 2467 2727 0 _1379_.A
rlabel metal2 2473 2753 2487 2767 0 _1379_.Y
rlabel metal1 2504 2642 2616 2658 0 _1380_.gnd
rlabel metal1 2504 2882 2616 2898 0 _1380_.vdd
rlabel metal2 2513 2733 2527 2747 0 _1380_.A
rlabel metal2 2573 2733 2587 2747 0 _1380_.Y
rlabel metal2 2553 2773 2567 2787 0 _1380_.B
rlabel metal1 2884 2642 3136 2658 0 _1566_.gnd
rlabel metal1 2884 2882 3136 2898 0 _1566_.vdd
rlabel metal2 2973 2733 2987 2747 0 _1566_.D
rlabel metal2 3013 2733 3027 2747 0 _1566_.CLK
rlabel metal2 3093 2733 3107 2747 0 _1566_.Q
rlabel metal1 2704 2642 2816 2658 0 _1382_.gnd
rlabel metal1 2704 2882 2816 2898 0 _1382_.vdd
rlabel metal2 2713 2733 2727 2747 0 _1382_.A
rlabel metal2 2733 2753 2747 2767 0 _1382_.B
rlabel metal2 2773 2753 2787 2767 0 _1382_.C
rlabel metal2 2753 2733 2767 2747 0 _1382_.Y
rlabel metal1 2804 2642 2896 2658 0 _1371_.gnd
rlabel metal1 2804 2882 2896 2898 0 _1371_.vdd
rlabel metal2 2813 2773 2827 2787 0 _1371_.A
rlabel metal2 2853 2773 2867 2787 0 _1371_.B
rlabel metal2 2833 2753 2847 2767 0 _1371_.Y
rlabel metal1 3124 2642 3376 2658 0 _1567_.gnd
rlabel metal1 3124 2882 3376 2898 0 _1567_.vdd
rlabel metal2 3213 2733 3227 2747 0 _1567_.D
rlabel metal2 3253 2733 3267 2747 0 _1567_.CLK
rlabel metal2 3333 2733 3347 2747 0 _1567_.Q
rlabel metal1 3424 2642 3516 2658 0 _1444_.gnd
rlabel metal1 3424 2882 3516 2898 0 _1444_.vdd
rlabel metal2 3453 2733 3467 2747 0 _1444_.B
rlabel metal2 3493 2733 3507 2747 0 _1444_.A
rlabel metal2 3473 2713 3487 2727 0 _1444_.Y
rlabel metal1 3364 2642 3436 2658 0 _1501_.gnd
rlabel metal1 3364 2882 3436 2898 0 _1501_.vdd
rlabel metal2 3413 2713 3427 2727 0 _1501_.A
rlabel metal2 3393 2753 3407 2767 0 _1501_.Y
rlabel metal1 3564 2642 3816 2658 0 _1598_.gnd
rlabel metal1 3564 2882 3816 2898 0 _1598_.vdd
rlabel metal2 3653 2733 3667 2747 0 _1598_.D
rlabel metal2 3693 2733 3707 2747 0 _1598_.CLK
rlabel metal2 3773 2733 3787 2747 0 _1598_.Q
rlabel metal1 3504 2642 3576 2658 0 _764_.gnd
rlabel metal1 3504 2882 3576 2898 0 _764_.vdd
rlabel metal2 3553 2753 3567 2767 0 _764_.A
rlabel metal2 3533 2733 3547 2747 0 _764_.Y
rlabel metal1 4004 2642 4116 2658 0 _767_.gnd
rlabel metal1 4004 2882 4116 2898 0 _767_.vdd
rlabel metal2 4013 2733 4027 2747 0 _767_.A
rlabel metal2 4033 2753 4047 2767 0 _767_.B
rlabel metal2 4073 2753 4087 2767 0 _767_.C
rlabel metal2 4053 2733 4067 2747 0 _767_.Y
rlabel metal1 3924 2642 4016 2658 0 _760_.gnd
rlabel metal1 3924 2882 4016 2898 0 _760_.vdd
rlabel metal2 3953 2733 3967 2747 0 _760_.B
rlabel metal2 3993 2733 4007 2747 0 _760_.A
rlabel metal2 3973 2713 3987 2727 0 _760_.Y
rlabel metal1 3804 2642 3936 2658 0 _776_.gnd
rlabel metal1 3804 2882 3936 2898 0 _776_.vdd
rlabel metal2 3913 2733 3927 2747 0 _776_.A
rlabel metal2 3893 2753 3907 2767 0 _776_.B
rlabel metal2 3833 2733 3847 2747 0 _776_.C
rlabel metal2 3853 2753 3867 2767 0 _776_.D
rlabel metal2 3873 2733 3887 2747 0 _776_.Y
rlabel metal1 4104 2642 4216 2658 0 _777_.gnd
rlabel metal1 4104 2882 4216 2898 0 _777_.vdd
rlabel metal2 4193 2733 4207 2747 0 _777_.A
rlabel metal2 4173 2753 4187 2767 0 _777_.B
rlabel metal2 4133 2753 4147 2767 0 _777_.C
rlabel metal2 4153 2733 4167 2747 0 _777_.Y
rlabel metal1 4204 2642 4296 2658 0 _774_.gnd
rlabel metal1 4204 2882 4296 2898 0 _774_.vdd
rlabel metal2 4253 2733 4267 2747 0 _774_.B
rlabel metal2 4213 2733 4227 2747 0 _774_.A
rlabel metal2 4233 2713 4247 2727 0 _774_.Y
rlabel metal1 4284 2642 4536 2658 0 _1577_.gnd
rlabel metal1 4284 2882 4536 2898 0 _1577_.vdd
rlabel metal2 4373 2733 4387 2747 0 _1577_.D
rlabel metal2 4413 2733 4427 2747 0 _1577_.CLK
rlabel metal2 4493 2733 4507 2747 0 _1577_.Q
rlabel metal1 4524 2642 4636 2658 0 _1485_.gnd
rlabel metal1 4524 2882 4636 2898 0 _1485_.vdd
rlabel metal2 4533 2733 4547 2747 0 _1485_.A
rlabel metal2 4553 2753 4567 2767 0 _1485_.B
rlabel metal2 4593 2753 4607 2767 0 _1485_.C
rlabel metal2 4573 2733 4587 2747 0 _1485_.Y
rlabel nsubstratencontact 4756 2888 4756 2888 0 FILL71250x39750.vdd
rlabel metal1 4744 2642 4776 2658 0 FILL71250x39750.gnd
rlabel nsubstratencontact 4736 2888 4736 2888 0 FILL70950x39750.vdd
rlabel metal1 4724 2642 4756 2658 0 FILL70950x39750.gnd
rlabel nsubstratencontact 4716 2888 4716 2888 0 FILL70650x39750.vdd
rlabel metal1 4704 2642 4736 2658 0 FILL70650x39750.gnd
rlabel metal1 4624 2642 4716 2658 0 _1484_.gnd
rlabel metal1 4624 2882 4716 2898 0 _1484_.vdd
rlabel metal2 4633 2773 4647 2787 0 _1484_.A
rlabel metal2 4673 2773 4687 2787 0 _1484_.B
rlabel metal2 4653 2753 4667 2767 0 _1484_.Y
rlabel metal1 4 3122 256 3138 0 _1596_.gnd
rlabel metal1 4 3362 256 3378 0 _1596_.vdd
rlabel metal2 93 3213 107 3227 0 _1596_.D
rlabel metal2 133 3213 147 3227 0 _1596_.CLK
rlabel metal2 213 3213 227 3227 0 _1596_.Q
rlabel metal1 224 3122 476 3138 0 _1527_.gnd
rlabel metal1 224 2882 476 2898 0 _1527_.vdd
rlabel metal2 373 3033 387 3047 0 _1527_.D
rlabel metal2 333 3033 347 3047 0 _1527_.CLK
rlabel metal2 253 3033 267 3047 0 _1527_.Q
rlabel metal1 244 3122 376 3138 0 _1161_.gnd
rlabel metal1 244 3362 376 3378 0 _1161_.vdd
rlabel metal2 353 3213 367 3227 0 _1161_.A
rlabel metal2 333 3233 347 3247 0 _1161_.B
rlabel metal2 273 3213 287 3227 0 _1161_.C
rlabel metal2 293 3233 307 3247 0 _1161_.D
rlabel metal2 313 3213 327 3227 0 _1161_.Y
rlabel metal1 4 3122 136 3138 0 _1158_.gnd
rlabel metal1 4 2882 136 2898 0 _1158_.vdd
rlabel metal2 113 3033 127 3047 0 _1158_.A
rlabel metal2 93 3013 107 3027 0 _1158_.B
rlabel metal2 33 3033 47 3047 0 _1158_.C
rlabel metal2 53 3013 67 3027 0 _1158_.D
rlabel metal2 73 3033 87 3047 0 _1158_.Y
rlabel metal1 124 3122 236 3138 0 _1157_.gnd
rlabel metal1 124 2882 236 2898 0 _1157_.vdd
rlabel metal2 213 3033 227 3047 0 _1157_.A
rlabel metal2 153 3033 167 3047 0 _1157_.Y
rlabel metal2 173 2993 187 3007 0 _1157_.B
rlabel metal1 444 3122 696 3138 0 _1529_.gnd
rlabel metal1 444 3362 696 3378 0 _1529_.vdd
rlabel metal2 593 3213 607 3227 0 _1529_.D
rlabel metal2 553 3213 567 3227 0 _1529_.CLK
rlabel metal2 473 3213 487 3227 0 _1529_.Q
rlabel metal1 464 3122 576 3138 0 _798_.gnd
rlabel metal1 464 2882 576 2898 0 _798_.vdd
rlabel metal2 473 3033 487 3047 0 _798_.A
rlabel metal2 493 3013 507 3027 0 _798_.B
rlabel metal2 533 3013 547 3027 0 _798_.C
rlabel metal2 513 3033 527 3047 0 _798_.Y
rlabel metal1 364 3122 456 3138 0 _1160_.gnd
rlabel metal1 364 3362 456 3378 0 _1160_.vdd
rlabel metal2 433 3253 447 3267 0 _1160_.A
rlabel metal2 393 3253 407 3267 0 _1160_.B
rlabel metal2 413 3233 427 3247 0 _1160_.Y
rlabel metal1 684 3122 796 3138 0 _802_.gnd
rlabel metal1 684 3362 796 3378 0 _802_.vdd
rlabel metal2 773 3213 787 3227 0 _802_.A
rlabel metal2 753 3233 767 3247 0 _802_.B
rlabel metal2 713 3233 727 3247 0 _802_.C
rlabel metal2 733 3213 747 3227 0 _802_.Y
rlabel metal1 644 3122 736 3138 0 _1520_.gnd
rlabel metal1 644 2882 736 2898 0 _1520_.vdd
rlabel metal2 713 2993 727 3007 0 _1520_.A
rlabel metal2 673 2993 687 3007 0 _1520_.B
rlabel metal2 693 3013 707 3027 0 _1520_.Y
rlabel metal1 564 3122 656 3138 0 _797_.gnd
rlabel metal1 564 2882 656 2898 0 _797_.vdd
rlabel metal2 573 2993 587 3007 0 _797_.A
rlabel metal2 613 2993 627 3007 0 _797_.B
rlabel metal2 593 3013 607 3027 0 _797_.Y
rlabel metal1 724 3122 816 3138 0 _1154_.gnd
rlabel metal1 724 2882 816 2898 0 _1154_.vdd
rlabel metal2 753 3033 767 3047 0 _1154_.B
rlabel metal2 793 3033 807 3047 0 _1154_.A
rlabel metal2 773 3053 787 3067 0 _1154_.Y
rlabel metal1 784 3122 916 3138 0 _1150_.gnd
rlabel metal1 784 3362 916 3378 0 _1150_.vdd
rlabel metal2 893 3213 907 3227 0 _1150_.A
rlabel metal2 873 3233 887 3247 0 _1150_.B
rlabel metal2 813 3213 827 3227 0 _1150_.C
rlabel metal2 833 3233 847 3247 0 _1150_.D
rlabel metal2 853 3213 867 3227 0 _1150_.Y
rlabel metal1 884 3122 996 3138 0 _1214_.gnd
rlabel metal1 884 2882 996 2898 0 _1214_.vdd
rlabel metal2 973 3033 987 3047 0 _1214_.A
rlabel metal2 953 3013 967 3027 0 _1214_.B
rlabel metal2 913 3013 927 3027 0 _1214_.C
rlabel metal2 933 3033 947 3047 0 _1214_.Y
rlabel metal1 984 3122 1096 3138 0 _1210_.gnd
rlabel metal1 984 2882 1096 2898 0 _1210_.vdd
rlabel metal2 1073 3033 1087 3047 0 _1210_.A
rlabel metal2 1053 3013 1067 3027 0 _1210_.B
rlabel metal2 1013 3013 1027 3027 0 _1210_.C
rlabel metal2 1033 3033 1047 3047 0 _1210_.Y
rlabel metal1 904 3122 996 3138 0 _1253_.gnd
rlabel metal1 904 3362 996 3378 0 _1253_.vdd
rlabel metal2 913 3253 927 3267 0 _1253_.A
rlabel metal2 953 3253 967 3267 0 _1253_.B
rlabel metal2 933 3233 947 3247 0 _1253_.Y
rlabel metal1 804 3122 896 3138 0 _1153_.gnd
rlabel metal1 804 2882 896 2898 0 _1153_.vdd
rlabel metal2 813 2993 827 3007 0 _1153_.A
rlabel metal2 853 2993 867 3007 0 _1153_.B
rlabel metal2 833 3013 847 3027 0 _1153_.Y
rlabel metal1 984 3122 1096 3138 0 _1149_.gnd
rlabel metal1 984 3362 1096 3378 0 _1149_.vdd
rlabel metal2 1073 3233 1087 3247 0 _1149_.A
rlabel metal2 1053 3253 1067 3267 0 _1149_.B
rlabel metal2 1033 3233 1047 3247 0 _1149_.C
rlabel metal2 1013 3253 1027 3267 0 _1149_.Y
rlabel metal1 1284 3122 1396 3138 0 _1247_.gnd
rlabel metal1 1284 3362 1396 3378 0 _1247_.vdd
rlabel metal2 1293 3213 1307 3227 0 _1247_.A
rlabel metal2 1313 3233 1327 3247 0 _1247_.B
rlabel metal2 1353 3233 1367 3247 0 _1247_.C
rlabel metal2 1333 3213 1347 3227 0 _1247_.Y
rlabel metal1 1164 3122 1276 3138 0 _1213_.gnd
rlabel metal1 1164 2882 1276 2898 0 _1213_.vdd
rlabel metal2 1253 3033 1267 3047 0 _1213_.A
rlabel metal2 1233 3013 1247 3027 0 _1213_.B
rlabel metal2 1193 3013 1207 3027 0 _1213_.C
rlabel metal2 1213 3033 1227 3047 0 _1213_.Y
rlabel metal1 1264 3122 1356 3138 0 _1212_.gnd
rlabel metal1 1264 2882 1356 2898 0 _1212_.vdd
rlabel metal2 1273 2993 1287 3007 0 _1212_.A
rlabel metal2 1313 2993 1327 3007 0 _1212_.B
rlabel metal2 1293 3013 1307 3027 0 _1212_.Y
rlabel metal1 1084 3122 1176 3138 0 _1206_.gnd
rlabel metal1 1084 2882 1176 2898 0 _1206_.vdd
rlabel metal2 1113 3033 1127 3047 0 _1206_.B
rlabel metal2 1153 3033 1167 3047 0 _1206_.A
rlabel metal2 1133 3053 1147 3067 0 _1206_.Y
rlabel metal1 1184 3122 1296 3138 0 _1211_.gnd
rlabel metal1 1184 3362 1296 3378 0 _1211_.vdd
rlabel metal2 1193 3233 1207 3247 0 _1211_.A
rlabel metal2 1213 3253 1227 3267 0 _1211_.B
rlabel metal2 1233 3233 1247 3247 0 _1211_.C
rlabel metal2 1253 3253 1267 3267 0 _1211_.Y
rlabel metal1 1084 3122 1196 3138 0 _1148_.gnd
rlabel metal1 1084 3362 1196 3378 0 _1148_.vdd
rlabel metal2 1173 3213 1187 3227 0 _1148_.A
rlabel metal2 1113 3213 1127 3227 0 _1148_.Y
rlabel metal2 1133 3253 1147 3267 0 _1148_.B
rlabel metal1 1564 3122 1656 3138 0 BUFX2_insert25.gnd
rlabel metal1 1564 2882 1656 2898 0 BUFX2_insert25.vdd
rlabel metal2 1573 3033 1587 3047 0 BUFX2_insert25.A
rlabel metal2 1613 3033 1627 3047 0 BUFX2_insert25.Y
rlabel metal1 1564 3122 1656 3138 0 _1257_.gnd
rlabel metal1 1564 3362 1656 3378 0 _1257_.vdd
rlabel metal2 1633 3253 1647 3267 0 _1257_.A
rlabel metal2 1593 3253 1607 3267 0 _1257_.B
rlabel metal2 1613 3233 1627 3247 0 _1257_.Y
rlabel metal1 1404 3122 1496 3138 0 _1250_.gnd
rlabel metal1 1404 2882 1496 2898 0 _1250_.vdd
rlabel metal2 1413 2993 1427 3007 0 _1250_.A
rlabel metal2 1453 2993 1467 3007 0 _1250_.B
rlabel metal2 1433 3013 1447 3027 0 _1250_.Y
rlabel metal1 1384 3122 1476 3138 0 _1209_.gnd
rlabel metal1 1384 3362 1476 3378 0 _1209_.vdd
rlabel metal2 1393 3253 1407 3267 0 _1209_.A
rlabel metal2 1433 3253 1447 3267 0 _1209_.B
rlabel metal2 1413 3233 1427 3247 0 _1209_.Y
rlabel metal1 1484 3122 1576 3138 0 _1207_.gnd
rlabel metal1 1484 2882 1576 2898 0 _1207_.vdd
rlabel metal2 1493 2993 1507 3007 0 _1207_.A
rlabel metal2 1533 2993 1547 3007 0 _1207_.B
rlabel metal2 1513 3013 1527 3027 0 _1207_.Y
rlabel metal1 1464 3122 1576 3138 0 _1255_.gnd
rlabel metal1 1464 3362 1576 3378 0 _1255_.vdd
rlabel metal2 1553 3193 1567 3207 0 _1255_.A
rlabel metal2 1533 3213 1547 3227 0 _1255_.B
rlabel metal2 1493 3233 1507 3247 0 _1255_.Y
rlabel metal1 1344 3122 1416 3138 0 _1146_.gnd
rlabel metal1 1344 2882 1416 2898 0 _1146_.vdd
rlabel metal2 1393 3013 1407 3027 0 _1146_.A
rlabel metal2 1373 3033 1387 3047 0 _1146_.Y
rlabel metal1 1644 3122 1756 3138 0 _1256_.gnd
rlabel metal1 1644 3362 1756 3378 0 _1256_.vdd
rlabel metal2 1653 3213 1667 3227 0 _1256_.A
rlabel metal2 1673 3233 1687 3247 0 _1256_.B
rlabel metal2 1713 3233 1727 3247 0 _1256_.C
rlabel metal2 1693 3213 1707 3227 0 _1256_.Y
rlabel metal1 1744 3122 1856 3138 0 _1254_.gnd
rlabel metal1 1744 3362 1856 3378 0 _1254_.vdd
rlabel metal2 1833 3213 1847 3227 0 _1254_.A
rlabel metal2 1813 3233 1827 3247 0 _1254_.B
rlabel metal2 1773 3233 1787 3247 0 _1254_.C
rlabel metal2 1793 3213 1807 3227 0 _1254_.Y
rlabel metal1 1644 3122 1756 3138 0 _1252_.gnd
rlabel metal1 1644 2882 1756 2898 0 _1252_.vdd
rlabel metal2 1653 3033 1667 3047 0 _1252_.A
rlabel metal2 1673 3013 1687 3027 0 _1252_.B
rlabel metal2 1713 3013 1727 3027 0 _1252_.C
rlabel metal2 1693 3033 1707 3047 0 _1252_.Y
rlabel metal1 1744 3122 1856 3138 0 _785_.gnd
rlabel metal1 1744 2882 1856 2898 0 _785_.vdd
rlabel metal2 1753 3033 1767 3047 0 _785_.A
rlabel metal2 1773 3013 1787 3027 0 _785_.B
rlabel metal2 1813 3013 1827 3027 0 _785_.C
rlabel metal2 1793 3033 1807 3047 0 _785_.Y
rlabel metal1 1844 3122 1936 3138 0 _1251_.gnd
rlabel metal1 1844 3362 1936 3378 0 _1251_.vdd
rlabel metal2 1853 3253 1867 3267 0 _1251_.A
rlabel metal2 1893 3253 1907 3267 0 _1251_.B
rlabel metal2 1873 3233 1887 3247 0 _1251_.Y
rlabel metal1 1844 3122 1936 3138 0 _1280_.gnd
rlabel metal1 1844 2882 1936 2898 0 _1280_.vdd
rlabel metal2 1893 3033 1907 3047 0 _1280_.B
rlabel metal2 1853 3033 1867 3047 0 _1280_.A
rlabel metal2 1873 3053 1887 3067 0 _1280_.Y
rlabel metal1 2084 3122 2196 3138 0 _1315_.gnd
rlabel metal1 2084 2882 2196 2898 0 _1315_.vdd
rlabel metal2 2093 3033 2107 3047 0 _1315_.A
rlabel metal2 2113 3013 2127 3027 0 _1315_.B
rlabel metal2 2153 3013 2167 3027 0 _1315_.C
rlabel metal2 2133 3033 2147 3047 0 _1315_.Y
rlabel metal1 2024 3122 2136 3138 0 _1279_.gnd
rlabel metal1 2024 3362 2136 3378 0 _1279_.vdd
rlabel metal2 2113 3213 2127 3227 0 _1279_.A
rlabel metal2 2093 3233 2107 3247 0 _1279_.B
rlabel metal2 2053 3233 2067 3247 0 _1279_.C
rlabel metal2 2073 3213 2087 3227 0 _1279_.Y
rlabel metal1 1924 3122 2036 3138 0 _1278_.gnd
rlabel metal1 1924 3362 2036 3378 0 _1278_.vdd
rlabel metal2 1933 3213 1947 3227 0 _1278_.A
rlabel metal2 1953 3233 1967 3247 0 _1278_.B
rlabel metal2 1993 3233 2007 3247 0 _1278_.C
rlabel metal2 1973 3213 1987 3227 0 _1278_.Y
rlabel metal1 1924 3122 2036 3138 0 _1271_.gnd
rlabel metal1 1924 2882 2036 2898 0 _1271_.vdd
rlabel metal2 1933 3013 1947 3027 0 _1271_.A
rlabel metal2 1953 3053 1967 3067 0 _1271_.B
rlabel metal2 1973 3013 1987 3027 0 _1271_.C
rlabel metal2 1993 3033 2007 3047 0 _1271_.Y
rlabel metal1 2024 3122 2096 3138 0 _1305_.gnd
rlabel metal1 2024 2882 2096 2898 0 _1305_.vdd
rlabel metal2 2033 3053 2047 3067 0 _1305_.A
rlabel metal2 2053 3013 2067 3027 0 _1305_.Y
rlabel metal1 2124 3122 2196 3138 0 _1208_.gnd
rlabel metal1 2124 3362 2196 3378 0 _1208_.vdd
rlabel metal2 2133 3193 2147 3207 0 _1208_.A
rlabel metal2 2153 3233 2167 3247 0 _1208_.Y
rlabel metal1 2184 3122 2296 3138 0 _1306_.gnd
rlabel metal1 2184 3362 2296 3378 0 _1306_.vdd
rlabel metal2 2193 3213 2207 3227 0 _1306_.A
rlabel metal2 2213 3233 2227 3247 0 _1306_.B
rlabel metal2 2253 3233 2267 3247 0 _1306_.C
rlabel metal2 2233 3213 2247 3227 0 _1306_.Y
rlabel metal1 2344 3122 2456 3138 0 _791_.gnd
rlabel metal1 2344 2882 2456 2898 0 _791_.vdd
rlabel metal2 2353 3033 2367 3047 0 _791_.A
rlabel metal2 2373 3013 2387 3027 0 _791_.B
rlabel metal2 2413 3013 2427 3027 0 _791_.C
rlabel metal2 2393 3033 2407 3047 0 _791_.Y
rlabel metal1 2344 3122 2436 3138 0 _1307_.gnd
rlabel metal1 2344 3362 2436 3378 0 _1307_.vdd
rlabel metal2 2353 3253 2367 3267 0 _1307_.A
rlabel metal2 2393 3253 2407 3267 0 _1307_.B
rlabel metal2 2373 3233 2387 3247 0 _1307_.Y
rlabel metal1 2264 3122 2356 3138 0 _790_.gnd
rlabel metal1 2264 2882 2356 2898 0 _790_.vdd
rlabel metal2 2333 2993 2347 3007 0 _790_.A
rlabel metal2 2293 2993 2307 3007 0 _790_.B
rlabel metal2 2313 3013 2327 3027 0 _790_.Y
rlabel metal1 2184 3122 2276 3138 0 _1316_.gnd
rlabel metal1 2184 2882 2276 2898 0 _1316_.vdd
rlabel metal2 2233 3033 2247 3047 0 _1316_.B
rlabel metal2 2193 3033 2207 3047 0 _1316_.A
rlabel metal2 2213 3053 2227 3067 0 _1316_.Y
rlabel metal1 2284 3122 2356 3138 0 _1314_.gnd
rlabel metal1 2284 3362 2356 3378 0 _1314_.vdd
rlabel metal2 2333 3193 2347 3207 0 _1314_.A
rlabel metal2 2313 3233 2327 3247 0 _1314_.Y
rlabel metal1 2664 3122 2756 3138 0 BUFX2_insert26.gnd
rlabel metal1 2664 3362 2756 3378 0 BUFX2_insert26.vdd
rlabel metal2 2673 3213 2687 3227 0 BUFX2_insert26.A
rlabel metal2 2713 3213 2727 3227 0 BUFX2_insert26.Y
rlabel metal1 2604 3122 2696 3138 0 BUFX2_insert1.gnd
rlabel metal1 2604 2882 2696 2898 0 BUFX2_insert1.vdd
rlabel metal2 2613 3033 2627 3047 0 BUFX2_insert1.A
rlabel metal2 2653 3033 2667 3047 0 BUFX2_insert1.Y
rlabel metal1 2424 3122 2676 3138 0 _1536_.gnd
rlabel metal1 2424 3362 2676 3378 0 _1536_.vdd
rlabel metal2 2573 3213 2587 3227 0 _1536_.D
rlabel metal2 2533 3213 2547 3227 0 _1536_.CLK
rlabel metal2 2453 3213 2467 3227 0 _1536_.Q
rlabel metal1 2504 3122 2616 3138 0 _823_.gnd
rlabel metal1 2504 2882 2616 2898 0 _823_.vdd
rlabel metal2 2513 3033 2527 3047 0 _823_.A
rlabel metal2 2533 3013 2547 3027 0 _823_.B
rlabel metal2 2573 3013 2587 3027 0 _823_.C
rlabel metal2 2553 3033 2567 3047 0 _823_.Y
rlabel metal1 2444 3122 2516 3138 0 _821_.gnd
rlabel metal1 2444 2882 2516 2898 0 _821_.vdd
rlabel metal2 2453 3053 2467 3067 0 _821_.A
rlabel metal2 2473 3013 2487 3027 0 _821_.Y
rlabel metal1 2764 3122 3016 3138 0 _1590_.gnd
rlabel metal1 2764 2882 3016 2898 0 _1590_.vdd
rlabel metal2 2853 3033 2867 3047 0 _1590_.D
rlabel metal2 2893 3033 2907 3047 0 _1590_.CLK
rlabel metal2 2973 3033 2987 3047 0 _1590_.Q
rlabel metal1 2744 3122 2996 3138 0 _1586_.gnd
rlabel metal1 2744 3362 2996 3378 0 _1586_.vdd
rlabel metal2 2893 3213 2907 3227 0 _1586_.D
rlabel metal2 2853 3213 2867 3227 0 _1586_.CLK
rlabel metal2 2773 3213 2787 3227 0 _1586_.Q
rlabel metal1 2684 3122 2776 3138 0 _822_.gnd
rlabel metal1 2684 2882 2776 2898 0 _822_.vdd
rlabel metal2 2693 2993 2707 3007 0 _822_.A
rlabel metal2 2733 2993 2747 3007 0 _822_.B
rlabel metal2 2713 3013 2727 3027 0 _822_.Y
rlabel metal1 3084 3122 3196 3138 0 _1509_.gnd
rlabel metal1 3084 3362 3196 3378 0 _1509_.vdd
rlabel metal2 3173 3213 3187 3227 0 _1509_.A
rlabel metal2 3153 3233 3167 3247 0 _1509_.B
rlabel metal2 3113 3233 3127 3247 0 _1509_.C
rlabel metal2 3133 3213 3147 3227 0 _1509_.Y
rlabel metal1 2984 3122 3096 3138 0 _1508_.gnd
rlabel metal1 2984 3362 3096 3378 0 _1508_.vdd
rlabel metal2 3073 3213 3087 3227 0 _1508_.A
rlabel metal2 3053 3233 3067 3247 0 _1508_.B
rlabel metal2 3013 3233 3027 3247 0 _1508_.C
rlabel metal2 3033 3213 3047 3227 0 _1508_.Y
rlabel metal1 3184 3122 3296 3138 0 _1506_.gnd
rlabel metal1 3184 3362 3296 3378 0 _1506_.vdd
rlabel metal2 3193 3213 3207 3227 0 _1506_.A
rlabel metal2 3213 3233 3227 3247 0 _1506_.B
rlabel metal2 3253 3233 3267 3247 0 _1506_.C
rlabel metal2 3233 3213 3247 3227 0 _1506_.Y
rlabel metal1 3084 3122 3196 3138 0 _1515_.gnd
rlabel metal1 3084 2882 3196 2898 0 _1515_.vdd
rlabel metal2 3173 3013 3187 3027 0 _1515_.A
rlabel metal2 3153 3053 3167 3067 0 _1515_.B
rlabel metal2 3133 3013 3147 3027 0 _1515_.C
rlabel metal2 3113 3033 3127 3047 0 _1515_.Y
rlabel metal1 3184 3122 3276 3138 0 _1514_.gnd
rlabel metal1 3184 2882 3276 2898 0 _1514_.vdd
rlabel metal2 3233 3033 3247 3047 0 _1514_.B
rlabel metal2 3193 3033 3207 3047 0 _1514_.A
rlabel metal2 3213 3053 3227 3067 0 _1514_.Y
rlabel metal1 3004 3122 3096 3138 0 _765_.gnd
rlabel metal1 3004 2882 3096 2898 0 _765_.vdd
rlabel metal2 3033 3033 3047 3047 0 _765_.B
rlabel metal2 3073 3033 3087 3047 0 _765_.A
rlabel metal2 3053 3053 3067 3067 0 _765_.Y
rlabel metal1 3264 3122 3516 3138 0 _1568_.gnd
rlabel metal1 3264 2882 3516 2898 0 _1568_.vdd
rlabel metal2 3353 3033 3367 3047 0 _1568_.D
rlabel metal2 3393 3033 3407 3047 0 _1568_.CLK
rlabel metal2 3473 3033 3487 3047 0 _1568_.Q
rlabel metal1 3284 3122 3396 3138 0 _1507_.gnd
rlabel metal1 3284 3362 3396 3378 0 _1507_.vdd
rlabel metal2 3373 3213 3387 3227 0 _1507_.A
rlabel metal2 3353 3233 3367 3247 0 _1507_.B
rlabel metal2 3313 3233 3327 3247 0 _1507_.C
rlabel metal2 3333 3213 3347 3227 0 _1507_.Y
rlabel metal1 3384 3122 3496 3138 0 _1407_.gnd
rlabel metal1 3384 3362 3496 3378 0 _1407_.vdd
rlabel metal2 3393 3213 3407 3227 0 _1407_.A
rlabel metal2 3413 3233 3427 3247 0 _1407_.B
rlabel metal2 3453 3233 3467 3247 0 _1407_.C
rlabel metal2 3433 3213 3447 3227 0 _1407_.Y
rlabel metal1 3504 3122 3756 3138 0 _1597_.gnd
rlabel metal1 3504 2882 3756 2898 0 _1597_.vdd
rlabel metal2 3593 3033 3607 3047 0 _1597_.D
rlabel metal2 3633 3033 3647 3047 0 _1597_.CLK
rlabel metal2 3713 3033 3727 3047 0 _1597_.Q
rlabel metal1 3484 3122 3576 3138 0 _1443_.gnd
rlabel metal1 3484 3362 3576 3378 0 _1443_.vdd
rlabel metal2 3493 3253 3507 3267 0 _1443_.A
rlabel metal2 3533 3253 3547 3267 0 _1443_.B
rlabel metal2 3513 3233 3527 3247 0 _1443_.Y
rlabel metal1 3644 3122 3736 3138 0 _1442_.gnd
rlabel metal1 3644 3362 3736 3378 0 _1442_.vdd
rlabel metal2 3653 3253 3667 3267 0 _1442_.A
rlabel metal2 3693 3253 3707 3267 0 _1442_.B
rlabel metal2 3673 3233 3687 3247 0 _1442_.Y
rlabel metal1 3564 3122 3656 3138 0 _1441_.gnd
rlabel metal1 3564 3362 3656 3378 0 _1441_.vdd
rlabel metal2 3573 3253 3587 3267 0 _1441_.A
rlabel metal2 3613 3253 3627 3267 0 _1441_.B
rlabel metal2 3593 3233 3607 3247 0 _1441_.Y
rlabel metal1 3724 3122 3816 3138 0 _1393_.gnd
rlabel metal1 3724 3362 3816 3378 0 _1393_.vdd
rlabel metal2 3733 3253 3747 3267 0 _1393_.A
rlabel metal2 3773 3253 3787 3267 0 _1393_.B
rlabel metal2 3753 3233 3767 3247 0 _1393_.Y
rlabel metal1 3804 3122 3896 3138 0 _1602_.gnd
rlabel metal1 3804 3362 3896 3378 0 _1602_.vdd
rlabel metal2 3813 3213 3827 3227 0 _1602_.A
rlabel metal2 3853 3213 3867 3227 0 _1602_.Y
rlabel metal1 3824 3122 3936 3138 0 _782_.gnd
rlabel metal1 3824 2882 3936 2898 0 _782_.vdd
rlabel metal2 3913 3033 3927 3047 0 _782_.A
rlabel metal2 3893 3013 3907 3027 0 _782_.B
rlabel metal2 3853 3013 3867 3027 0 _782_.C
rlabel metal2 3873 3033 3887 3047 0 _782_.Y
rlabel metal1 3924 3122 4036 3138 0 _780_.gnd
rlabel metal1 3924 2882 4036 2898 0 _780_.vdd
rlabel metal2 4013 3033 4027 3047 0 _780_.A
rlabel metal2 3993 3013 4007 3027 0 _780_.B
rlabel metal2 3953 3013 3967 3027 0 _780_.C
rlabel metal2 3973 3033 3987 3047 0 _780_.Y
rlabel metal1 3884 3122 3976 3138 0 _779_.gnd
rlabel metal1 3884 3362 3976 3378 0 _779_.vdd
rlabel metal2 3953 3253 3967 3267 0 _779_.A
rlabel metal2 3913 3253 3927 3267 0 _779_.B
rlabel metal2 3933 3233 3947 3247 0 _779_.Y
rlabel metal1 3964 3122 4056 3138 0 _1492_.gnd
rlabel metal1 3964 3362 4056 3378 0 _1492_.vdd
rlabel metal2 3993 3213 4007 3227 0 _1492_.B
rlabel metal2 4033 3213 4047 3227 0 _1492_.A
rlabel metal2 4013 3193 4027 3207 0 _1492_.Y
rlabel metal1 3744 3122 3836 3138 0 _762_.gnd
rlabel metal1 3744 2882 3836 2898 0 _762_.vdd
rlabel metal2 3793 3033 3807 3047 0 _762_.B
rlabel metal2 3753 3033 3767 3047 0 _762_.A
rlabel metal2 3773 3053 3787 3067 0 _762_.Y
rlabel metal1 4044 3122 4136 3138 0 _1606_.gnd
rlabel metal1 4044 3362 4136 3378 0 _1606_.vdd
rlabel metal2 4053 3213 4067 3227 0 _1606_.A
rlabel metal2 4093 3213 4107 3227 0 _1606_.Y
rlabel metal1 4124 3122 4236 3138 0 _775_.gnd
rlabel metal1 4124 2882 4236 2898 0 _775_.vdd
rlabel metal2 4133 3033 4147 3047 0 _775_.A
rlabel metal2 4153 3013 4167 3027 0 _775_.B
rlabel metal2 4193 3013 4207 3027 0 _775_.C
rlabel metal2 4173 3033 4187 3047 0 _775_.Y
rlabel metal1 4184 3122 4296 3138 0 _773_.gnd
rlabel metal1 4184 3362 4296 3378 0 _773_.vdd
rlabel metal2 4273 3213 4287 3227 0 _773_.A
rlabel metal2 4253 3233 4267 3247 0 _773_.B
rlabel metal2 4213 3233 4227 3247 0 _773_.C
rlabel metal2 4233 3213 4247 3227 0 _773_.Y
rlabel metal1 4024 3122 4136 3138 0 _763_.gnd
rlabel metal1 4024 2882 4136 2898 0 _763_.vdd
rlabel metal2 4033 3033 4047 3047 0 _763_.A
rlabel metal2 4053 3013 4067 3027 0 _763_.B
rlabel metal2 4093 3013 4107 3027 0 _763_.C
rlabel metal2 4073 3033 4087 3047 0 _763_.Y
rlabel metal1 4224 3122 4296 3138 0 _768_.gnd
rlabel metal1 4224 2882 4296 2898 0 _768_.vdd
rlabel metal2 4233 3053 4247 3067 0 _768_.A
rlabel metal2 4253 3013 4267 3027 0 _768_.Y
rlabel metal1 4124 3122 4196 3138 0 _761_.gnd
rlabel metal1 4124 3362 4196 3378 0 _761_.vdd
rlabel metal2 4173 3193 4187 3207 0 _761_.A
rlabel metal2 4153 3233 4167 3247 0 _761_.Y
rlabel metal1 4384 3122 4636 3138 0 _1599_.gnd
rlabel metal1 4384 2882 4636 2898 0 _1599_.vdd
rlabel metal2 4533 3033 4547 3047 0 _1599_.D
rlabel metal2 4493 3033 4507 3047 0 _1599_.CLK
rlabel metal2 4413 3033 4427 3047 0 _1599_.Q
rlabel metal1 4524 3122 4776 3138 0 _1578_.gnd
rlabel metal1 4524 3362 4776 3378 0 _1578_.vdd
rlabel metal2 4613 3213 4627 3227 0 _1578_.D
rlabel metal2 4653 3213 4667 3227 0 _1578_.CLK
rlabel metal2 4733 3213 4747 3227 0 _1578_.Q
rlabel metal1 4344 3122 4456 3138 0 _771_.gnd
rlabel metal1 4344 3362 4456 3378 0 _771_.vdd
rlabel metal2 4353 3213 4367 3227 0 _771_.A
rlabel metal2 4373 3233 4387 3247 0 _771_.B
rlabel metal2 4413 3233 4427 3247 0 _771_.C
rlabel metal2 4393 3213 4407 3227 0 _771_.Y
rlabel metal1 4444 3122 4536 3138 0 _770_.gnd
rlabel metal1 4444 3362 4536 3378 0 _770_.vdd
rlabel metal2 4513 3253 4527 3267 0 _770_.A
rlabel metal2 4473 3253 4487 3267 0 _770_.B
rlabel metal2 4493 3233 4507 3247 0 _770_.Y
rlabel metal1 4284 3122 4356 3138 0 _1454_.gnd
rlabel metal1 4284 3362 4356 3378 0 _1454_.vdd
rlabel metal2 4333 3193 4347 3207 0 _1454_.A
rlabel metal2 4313 3233 4327 3247 0 _1454_.Y
rlabel metal1 4284 3122 4396 3138 0 _1480_.gnd
rlabel metal1 4284 2882 4396 2898 0 _1480_.vdd
rlabel metal2 4293 3013 4307 3027 0 _1480_.A
rlabel metal2 4313 2993 4327 3007 0 _1480_.B
rlabel metal2 4333 3013 4347 3027 0 _1480_.C
rlabel metal2 4353 2993 4367 3007 0 _1480_.Y
rlabel nsubstratencontact 4764 2892 4764 2892 0 FILL71250x43350.vdd
rlabel metal1 4744 3122 4776 3138 0 FILL71250x43350.gnd
rlabel nsubstratencontact 4744 2892 4744 2892 0 FILL70950x43350.vdd
rlabel metal1 4724 3122 4756 3138 0 FILL70950x43350.gnd
rlabel metal1 4624 3122 4736 3138 0 _1488_.gnd
rlabel metal1 4624 2882 4736 2898 0 _1488_.vdd
rlabel metal2 4633 3033 4647 3047 0 _1488_.A
rlabel metal2 4653 3013 4667 3027 0 _1488_.B
rlabel metal2 4693 3013 4707 3027 0 _1488_.C
rlabel metal2 4673 3033 4687 3047 0 _1488_.Y
rlabel metal1 84 3602 336 3618 0 _1595_.gnd
rlabel metal1 84 3362 336 3378 0 _1595_.vdd
rlabel metal2 173 3513 187 3527 0 _1595_.D
rlabel metal2 213 3513 227 3527 0 _1595_.CLK
rlabel metal2 293 3513 307 3527 0 _1595_.Q
rlabel metal1 4 3602 96 3618 0 _1159_.gnd
rlabel metal1 4 3362 96 3378 0 _1159_.vdd
rlabel metal2 73 3473 87 3487 0 _1159_.A
rlabel metal2 33 3473 47 3487 0 _1159_.B
rlabel metal2 53 3493 67 3507 0 _1159_.Y
rlabel metal1 464 3602 576 3618 0 _1525_.gnd
rlabel metal1 464 3362 576 3378 0 _1525_.vdd
rlabel metal2 553 3513 567 3527 0 _1525_.A
rlabel metal2 533 3493 547 3507 0 _1525_.B
rlabel metal2 493 3493 507 3507 0 _1525_.C
rlabel metal2 513 3513 527 3527 0 _1525_.Y
rlabel metal1 384 3602 476 3618 0 _1524_.gnd
rlabel metal1 384 3362 476 3378 0 _1524_.vdd
rlabel metal2 453 3473 467 3487 0 _1524_.A
rlabel metal2 413 3473 427 3487 0 _1524_.B
rlabel metal2 433 3493 447 3507 0 _1524_.Y
rlabel metal1 324 3602 396 3618 0 _1166_.gnd
rlabel metal1 324 3362 396 3378 0 _1166_.vdd
rlabel metal2 373 3533 387 3547 0 _1166_.A
rlabel metal2 353 3493 367 3507 0 _1166_.Y
rlabel metal1 564 3602 676 3618 0 _1217_.gnd
rlabel metal1 564 3362 676 3378 0 _1217_.vdd
rlabel metal2 653 3513 667 3527 0 _1217_.A
rlabel metal2 633 3493 647 3507 0 _1217_.B
rlabel metal2 593 3493 607 3507 0 _1217_.C
rlabel metal2 613 3513 627 3527 0 _1217_.Y
rlabel metal1 664 3602 756 3618 0 _801_.gnd
rlabel metal1 664 3362 756 3378 0 _801_.vdd
rlabel metal2 673 3473 687 3487 0 _801_.A
rlabel metal2 713 3473 727 3487 0 _801_.B
rlabel metal2 693 3493 707 3507 0 _801_.Y
rlabel metal1 744 3602 876 3618 0 _1155_.gnd
rlabel metal1 744 3362 876 3378 0 _1155_.vdd
rlabel metal2 753 3513 767 3527 0 _1155_.A
rlabel metal2 773 3493 787 3507 0 _1155_.B
rlabel metal2 833 3513 847 3527 0 _1155_.C
rlabel metal2 793 3513 807 3527 0 _1155_.Y
rlabel metal2 813 3493 827 3507 0 _1155_.D
rlabel metal1 1024 3602 1136 3618 0 _1202_.gnd
rlabel metal1 1024 3362 1136 3378 0 _1202_.vdd
rlabel metal2 1033 3493 1047 3507 0 _1202_.A
rlabel metal2 1053 3533 1067 3547 0 _1202_.B
rlabel metal2 1073 3493 1087 3507 0 _1202_.C
rlabel metal2 1093 3513 1107 3527 0 _1202_.Y
rlabel metal1 864 3602 936 3618 0 _1151_.gnd
rlabel metal1 864 3362 936 3378 0 _1151_.vdd
rlabel metal2 873 3533 887 3547 0 _1151_.A
rlabel metal2 893 3493 907 3507 0 _1151_.Y
rlabel metal1 924 3602 1036 3618 0 _1152_.gnd
rlabel metal1 924 3362 1036 3378 0 _1152_.vdd
rlabel metal2 1013 3493 1027 3507 0 _1152_.A
rlabel metal2 993 3473 1007 3487 0 _1152_.B
rlabel metal2 973 3493 987 3507 0 _1152_.C
rlabel metal2 953 3473 967 3487 0 _1152_.Y
rlabel metal1 1204 3602 1296 3618 0 _1522_.gnd
rlabel metal1 1204 3362 1296 3378 0 _1522_.vdd
rlabel metal2 1213 3473 1227 3487 0 _1522_.A
rlabel metal2 1253 3473 1267 3487 0 _1522_.B
rlabel metal2 1233 3493 1247 3507 0 _1522_.Y
rlabel metal1 1284 3602 1376 3618 0 _799_.gnd
rlabel metal1 1284 3362 1376 3378 0 _799_.vdd
rlabel metal2 1293 3473 1307 3487 0 _799_.A
rlabel metal2 1333 3473 1347 3487 0 _799_.B
rlabel metal2 1313 3493 1327 3507 0 _799_.Y
rlabel metal1 1124 3602 1216 3618 0 _1147_.gnd
rlabel metal1 1124 3362 1216 3378 0 _1147_.vdd
rlabel metal2 1173 3513 1187 3527 0 _1147_.B
rlabel metal2 1133 3513 1147 3527 0 _1147_.A
rlabel metal2 1153 3533 1167 3547 0 _1147_.Y
rlabel metal1 1464 3602 1716 3618 0 _1528_.gnd
rlabel metal1 1464 3362 1716 3378 0 _1528_.vdd
rlabel metal2 1553 3513 1567 3527 0 _1528_.D
rlabel metal2 1593 3513 1607 3527 0 _1528_.CLK
rlabel metal2 1673 3513 1687 3527 0 _1528_.Q
rlabel metal1 1364 3602 1476 3618 0 _800_.gnd
rlabel metal1 1364 3362 1476 3378 0 _800_.vdd
rlabel metal2 1373 3513 1387 3527 0 _800_.A
rlabel metal2 1393 3493 1407 3507 0 _800_.B
rlabel metal2 1433 3493 1447 3507 0 _800_.C
rlabel metal2 1413 3513 1427 3527 0 _800_.Y
rlabel metal1 1784 3602 1896 3618 0 _794_.gnd
rlabel metal1 1784 3362 1896 3378 0 _794_.vdd
rlabel metal2 1793 3513 1807 3527 0 _794_.A
rlabel metal2 1813 3493 1827 3507 0 _794_.B
rlabel metal2 1853 3493 1867 3507 0 _794_.C
rlabel metal2 1833 3513 1847 3527 0 _794_.Y
rlabel metal1 1704 3602 1796 3618 0 _793_.gnd
rlabel metal1 1704 3362 1796 3378 0 _793_.vdd
rlabel metal2 1773 3473 1787 3487 0 _793_.A
rlabel metal2 1733 3473 1747 3487 0 _793_.B
rlabel metal2 1753 3493 1767 3507 0 _793_.Y
rlabel metal1 1944 3602 2036 3618 0 _1284_.gnd
rlabel metal1 1944 3362 2036 3378 0 _1284_.vdd
rlabel metal2 2013 3473 2027 3487 0 _1284_.A
rlabel metal2 1973 3473 1987 3487 0 _1284_.B
rlabel metal2 1993 3493 2007 3507 0 _1284_.Y
rlabel metal1 2124 3602 2216 3618 0 _1281_.gnd
rlabel metal1 2124 3362 2216 3378 0 _1281_.vdd
rlabel metal2 2133 3473 2147 3487 0 _1281_.A
rlabel metal2 2173 3473 2187 3487 0 _1281_.B
rlabel metal2 2153 3493 2167 3507 0 _1281_.Y
rlabel metal1 2024 3602 2136 3618 0 _1282_.gnd
rlabel metal1 2024 3362 2136 3378 0 _1282_.vdd
rlabel metal2 2113 3513 2127 3527 0 _1282_.A
rlabel metal2 2053 3513 2067 3527 0 _1282_.Y
rlabel metal2 2073 3473 2087 3487 0 _1282_.B
rlabel metal1 1884 3602 1956 3618 0 _789_.gnd
rlabel metal1 1884 3362 1956 3378 0 _789_.vdd
rlabel metal2 1893 3493 1907 3507 0 _789_.A
rlabel metal2 1913 3513 1927 3527 0 _789_.Y
rlabel metal1 2304 3602 2376 3618 0 _1303_.gnd
rlabel metal1 2304 3362 2376 3378 0 _1303_.vdd
rlabel metal2 2313 3533 2327 3547 0 _1303_.A
rlabel metal2 2333 3493 2347 3507 0 _1303_.Y
rlabel metal1 2364 3602 2436 3618 0 _824_.gnd
rlabel metal1 2364 3362 2436 3378 0 _824_.vdd
rlabel metal2 2373 3533 2387 3547 0 _824_.A
rlabel metal2 2393 3493 2407 3507 0 _824_.Y
rlabel metal1 2204 3602 2316 3618 0 _1304_.gnd
rlabel metal1 2204 3362 2316 3378 0 _1304_.vdd
rlabel metal2 2213 3493 2227 3507 0 _1304_.A
rlabel metal2 2233 3473 2247 3487 0 _1304_.B
rlabel metal2 2253 3493 2267 3507 0 _1304_.C
rlabel metal2 2273 3473 2287 3487 0 _1304_.Y
rlabel metal1 2424 3602 2676 3618 0 _1537_.gnd
rlabel metal1 2424 3362 2676 3378 0 _1537_.vdd
rlabel metal2 2573 3513 2587 3527 0 _1537_.D
rlabel metal2 2533 3513 2547 3527 0 _1537_.CLK
rlabel metal2 2453 3513 2467 3527 0 _1537_.Q
rlabel metal1 2664 3602 2776 3618 0 _826_.gnd
rlabel metal1 2664 3362 2776 3378 0 _826_.vdd
rlabel metal2 2673 3513 2687 3527 0 _826_.A
rlabel metal2 2693 3493 2707 3507 0 _826_.B
rlabel metal2 2733 3493 2747 3507 0 _826_.C
rlabel metal2 2713 3513 2727 3527 0 _826_.Y
rlabel metal1 2764 3602 2856 3618 0 BUFX2_insert3.gnd
rlabel metal1 2764 3362 2856 3378 0 BUFX2_insert3.vdd
rlabel metal2 2773 3513 2787 3527 0 BUFX2_insert3.A
rlabel metal2 2813 3513 2827 3527 0 BUFX2_insert3.Y
rlabel metal1 2924 3602 3176 3618 0 _1587_.gnd
rlabel metal1 2924 3362 3176 3378 0 _1587_.vdd
rlabel metal2 3073 3513 3087 3527 0 _1587_.D
rlabel metal2 3033 3513 3047 3527 0 _1587_.CLK
rlabel metal2 2953 3513 2967 3527 0 _1587_.Q
rlabel metal1 2844 3602 2936 3618 0 _825_.gnd
rlabel metal1 2844 3362 2936 3378 0 _825_.vdd
rlabel metal2 2853 3473 2867 3487 0 _825_.A
rlabel metal2 2893 3473 2907 3487 0 _825_.B
rlabel metal2 2873 3493 2887 3507 0 _825_.Y
rlabel metal1 3164 3602 3276 3618 0 _1406_.gnd
rlabel metal1 3164 3362 3276 3378 0 _1406_.vdd
rlabel metal2 3253 3513 3267 3527 0 _1406_.A
rlabel metal2 3233 3493 3247 3507 0 _1406_.B
rlabel metal2 3193 3493 3207 3507 0 _1406_.C
rlabel metal2 3213 3513 3227 3527 0 _1406_.Y
rlabel metal1 3464 3602 3556 3618 0 _1440_.gnd
rlabel metal1 3464 3362 3556 3378 0 _1440_.vdd
rlabel metal2 3493 3513 3507 3527 0 _1440_.B
rlabel metal2 3533 3513 3547 3527 0 _1440_.A
rlabel metal2 3513 3533 3527 3547 0 _1440_.Y
rlabel metal1 3324 3602 3416 3618 0 _1404_.gnd
rlabel metal1 3324 3362 3416 3378 0 _1404_.vdd
rlabel metal2 3373 3513 3387 3527 0 _1404_.B
rlabel metal2 3333 3513 3347 3527 0 _1404_.A
rlabel metal2 3353 3533 3367 3547 0 _1404_.Y
rlabel metal1 3264 3602 3336 3618 0 _1405_.gnd
rlabel metal1 3264 3362 3336 3378 0 _1405_.vdd
rlabel metal2 3313 3533 3327 3547 0 _1405_.A
rlabel metal2 3293 3493 3307 3507 0 _1405_.Y
rlabel metal1 3404 3602 3476 3618 0 _1400_.gnd
rlabel metal1 3404 3362 3476 3378 0 _1400_.vdd
rlabel metal2 3413 3533 3427 3547 0 _1400_.A
rlabel metal2 3433 3493 3447 3507 0 _1400_.Y
rlabel metal1 3544 3602 3656 3618 0 _1436_.gnd
rlabel metal1 3544 3362 3656 3378 0 _1436_.vdd
rlabel metal2 3553 3493 3567 3507 0 _1436_.A
rlabel metal2 3573 3533 3587 3547 0 _1436_.B
rlabel metal2 3593 3493 3607 3507 0 _1436_.C
rlabel metal2 3613 3513 3627 3527 0 _1436_.Y
rlabel metal1 3644 3602 3756 3618 0 _1435_.gnd
rlabel metal1 3644 3362 3756 3378 0 _1435_.vdd
rlabel metal2 3653 3533 3667 3547 0 _1435_.A
rlabel metal2 3673 3513 3687 3527 0 _1435_.B
rlabel metal2 3713 3493 3727 3507 0 _1435_.Y
rlabel metal1 3944 3602 4196 3618 0 _1571_.gnd
rlabel metal1 3944 3362 4196 3378 0 _1571_.vdd
rlabel metal2 4093 3513 4107 3527 0 _1571_.D
rlabel metal2 4053 3513 4067 3527 0 _1571_.CLK
rlabel metal2 3973 3513 3987 3527 0 _1571_.Q
rlabel metal1 3864 3602 3956 3618 0 _1416_.gnd
rlabel metal1 3864 3362 3956 3378 0 _1416_.vdd
rlabel metal2 3933 3473 3947 3487 0 _1416_.A
rlabel metal2 3893 3473 3907 3487 0 _1416_.B
rlabel metal2 3913 3493 3927 3507 0 _1416_.Y
rlabel metal1 3744 3602 3876 3618 0 _1437_.gnd
rlabel metal1 3744 3362 3876 3378 0 _1437_.vdd
rlabel metal2 3853 3513 3867 3527 0 _1437_.A
rlabel metal2 3833 3493 3847 3507 0 _1437_.B
rlabel metal2 3773 3513 3787 3527 0 _1437_.C
rlabel metal2 3793 3493 3807 3507 0 _1437_.D
rlabel metal2 3813 3513 3827 3527 0 _1437_.Y
rlabel metal1 4184 3602 4436 3618 0 _1600_.gnd
rlabel metal1 4184 3362 4436 3378 0 _1600_.vdd
rlabel metal2 4333 3513 4347 3527 0 _1600_.D
rlabel metal2 4293 3513 4307 3527 0 _1600_.CLK
rlabel metal2 4213 3513 4227 3527 0 _1600_.Q
rlabel metal1 4424 3602 4636 3618 0 CLKBUF1_insert9.gnd
rlabel metal1 4424 3362 4636 3378 0 CLKBUF1_insert9.vdd
rlabel metal2 4593 3493 4607 3507 0 CLKBUF1_insert9.A
rlabel metal2 4453 3493 4467 3507 0 CLKBUF1_insert9.Y
rlabel nsubstratencontact 4764 3372 4764 3372 0 FILL71250x50550.vdd
rlabel metal1 4744 3602 4776 3618 0 FILL71250x50550.gnd
rlabel nsubstratencontact 4744 3372 4744 3372 0 FILL70950x50550.vdd
rlabel metal1 4724 3602 4756 3618 0 FILL70950x50550.gnd
rlabel metal1 4624 3602 4736 3618 0 _844_.gnd
rlabel metal1 4624 3362 4736 3378 0 _844_.vdd
rlabel metal2 4633 3513 4647 3527 0 _844_.A
rlabel metal2 4653 3493 4667 3507 0 _844_.B
rlabel metal2 4693 3493 4707 3507 0 _844_.C
rlabel metal2 4673 3513 4687 3527 0 _844_.Y
rlabel metal1 84 3602 196 3618 0 _1163_.gnd
rlabel metal1 84 3842 196 3858 0 _1163_.vdd
rlabel metal2 93 3693 107 3707 0 _1163_.A
rlabel metal2 113 3713 127 3727 0 _1163_.B
rlabel metal2 153 3713 167 3727 0 _1163_.C
rlabel metal2 133 3693 147 3707 0 _1163_.Y
rlabel metal1 244 3602 356 3618 0 _1167_.gnd
rlabel metal1 244 3842 356 3858 0 _1167_.vdd
rlabel metal2 333 3713 347 3727 0 _1167_.A
rlabel metal2 313 3673 327 3687 0 _1167_.B
rlabel metal2 293 3713 307 3727 0 _1167_.C
rlabel metal2 273 3693 287 3707 0 _1167_.Y
rlabel metal1 4 3602 96 3618 0 _1164_.gnd
rlabel metal1 4 3842 96 3858 0 _1164_.vdd
rlabel metal2 33 3693 47 3707 0 _1164_.B
rlabel metal2 73 3693 87 3707 0 _1164_.A
rlabel metal2 53 3673 67 3687 0 _1164_.Y
rlabel metal1 184 3602 256 3618 0 _1162_.gnd
rlabel metal1 184 3842 256 3858 0 _1162_.vdd
rlabel metal2 233 3673 247 3687 0 _1162_.A
rlabel metal2 213 3713 227 3727 0 _1162_.Y
rlabel metal1 524 3602 616 3618 0 _1249_.gnd
rlabel metal1 524 3842 616 3858 0 _1249_.vdd
rlabel metal2 593 3733 607 3747 0 _1249_.A
rlabel metal2 553 3733 567 3747 0 _1249_.B
rlabel metal2 573 3713 587 3727 0 _1249_.Y
rlabel metal1 444 3602 536 3618 0 _1156_.gnd
rlabel metal1 444 3842 536 3858 0 _1156_.vdd
rlabel metal2 513 3733 527 3747 0 _1156_.A
rlabel metal2 473 3733 487 3747 0 _1156_.B
rlabel metal2 493 3713 507 3727 0 _1156_.Y
rlabel metal1 344 3602 456 3618 0 _1170_.gnd
rlabel metal1 344 3842 456 3858 0 _1170_.vdd
rlabel metal2 433 3693 447 3707 0 _1170_.A
rlabel metal2 373 3693 387 3707 0 _1170_.Y
rlabel metal2 393 3733 407 3747 0 _1170_.B
rlabel metal1 664 3602 776 3618 0 _1216_.gnd
rlabel metal1 664 3842 776 3858 0 _1216_.vdd
rlabel metal2 673 3693 687 3707 0 _1216_.A
rlabel metal2 693 3713 707 3727 0 _1216_.B
rlabel metal2 733 3713 747 3727 0 _1216_.C
rlabel metal2 713 3693 727 3707 0 _1216_.Y
rlabel metal1 764 3602 856 3618 0 _1215_.gnd
rlabel metal1 764 3842 856 3858 0 _1215_.vdd
rlabel metal2 773 3733 787 3747 0 _1215_.A
rlabel metal2 813 3733 827 3747 0 _1215_.B
rlabel metal2 793 3713 807 3727 0 _1215_.Y
rlabel metal1 604 3602 676 3618 0 _1218_.gnd
rlabel metal1 604 3842 676 3858 0 _1218_.vdd
rlabel metal2 613 3673 627 3687 0 _1218_.A
rlabel metal2 633 3713 647 3727 0 _1218_.Y
rlabel metal1 944 3602 1056 3618 0 _1223_.gnd
rlabel metal1 944 3842 1056 3858 0 _1223_.vdd
rlabel metal2 953 3713 967 3727 0 _1223_.A
rlabel metal2 973 3673 987 3687 0 _1223_.B
rlabel metal2 993 3713 1007 3727 0 _1223_.C
rlabel metal2 1013 3693 1027 3707 0 _1223_.Y
rlabel metal1 1044 3602 1156 3618 0 _1259_.gnd
rlabel metal1 1044 3842 1156 3858 0 _1259_.vdd
rlabel metal2 1053 3713 1067 3727 0 _1259_.A
rlabel metal2 1073 3733 1087 3747 0 _1259_.B
rlabel metal2 1093 3713 1107 3727 0 _1259_.C
rlabel metal2 1113 3733 1127 3747 0 _1259_.Y
rlabel metal1 844 3602 956 3618 0 _1219_.gnd
rlabel metal1 844 3842 956 3858 0 _1219_.vdd
rlabel metal2 933 3713 947 3727 0 _1219_.A
rlabel metal2 913 3733 927 3747 0 _1219_.B
rlabel metal2 893 3713 907 3727 0 _1219_.C
rlabel metal2 873 3733 887 3747 0 _1219_.Y
rlabel metal1 1144 3602 1256 3618 0 _1258_.gnd
rlabel metal1 1144 3842 1256 3858 0 _1258_.vdd
rlabel metal2 1153 3713 1167 3727 0 _1258_.A
rlabel metal2 1173 3673 1187 3687 0 _1258_.B
rlabel metal2 1193 3713 1207 3727 0 _1258_.C
rlabel metal2 1213 3693 1227 3707 0 _1258_.Y
rlabel metal1 1244 3602 1316 3618 0 _1262_.gnd
rlabel metal1 1244 3842 1316 3858 0 _1262_.vdd
rlabel metal2 1253 3673 1267 3687 0 _1262_.A
rlabel metal2 1273 3713 1287 3727 0 _1262_.Y
rlabel metal1 1304 3602 1416 3618 0 _1263_.gnd
rlabel metal1 1304 3842 1416 3858 0 _1263_.vdd
rlabel metal2 1393 3713 1407 3727 0 _1263_.A
rlabel metal2 1373 3733 1387 3747 0 _1263_.B
rlabel metal2 1353 3713 1367 3727 0 _1263_.C
rlabel metal2 1333 3733 1347 3747 0 _1263_.Y
rlabel metal1 1464 3602 1576 3618 0 _1261_.gnd
rlabel metal1 1464 3842 1576 3858 0 _1261_.vdd
rlabel metal2 1553 3693 1567 3707 0 _1261_.A
rlabel metal2 1533 3713 1547 3727 0 _1261_.B
rlabel metal2 1493 3713 1507 3727 0 _1261_.C
rlabel metal2 1513 3693 1527 3707 0 _1261_.Y
rlabel metal1 1564 3602 1636 3618 0 _1260_.gnd
rlabel metal1 1564 3842 1636 3858 0 _1260_.vdd
rlabel metal2 1613 3673 1627 3687 0 _1260_.A
rlabel metal2 1593 3713 1607 3727 0 _1260_.Y
rlabel metal1 1404 3602 1476 3618 0 _1248_.gnd
rlabel metal1 1404 3842 1476 3858 0 _1248_.vdd
rlabel metal2 1453 3673 1467 3687 0 _1248_.A
rlabel metal2 1433 3713 1447 3727 0 _1248_.Y
rlabel metal1 1804 3602 1916 3618 0 _1302_.gnd
rlabel metal1 1804 3842 1916 3858 0 _1302_.vdd
rlabel metal2 1893 3713 1907 3727 0 _1302_.A
rlabel metal2 1873 3673 1887 3687 0 _1302_.B
rlabel metal2 1853 3713 1867 3727 0 _1302_.C
rlabel metal2 1833 3693 1847 3707 0 _1302_.Y
rlabel metal1 1624 3602 1736 3618 0 _1277_.gnd
rlabel metal1 1624 3842 1736 3858 0 _1277_.vdd
rlabel metal2 1633 3713 1647 3727 0 _1277_.A
rlabel metal2 1653 3673 1667 3687 0 _1277_.B
rlabel metal2 1673 3713 1687 3727 0 _1277_.C
rlabel metal2 1693 3693 1707 3707 0 _1277_.Y
rlabel metal1 1724 3602 1816 3618 0 _1286_.gnd
rlabel metal1 1724 3842 1816 3858 0 _1286_.vdd
rlabel metal2 1773 3693 1787 3707 0 _1286_.B
rlabel metal2 1733 3693 1747 3707 0 _1286_.A
rlabel metal2 1753 3673 1767 3687 0 _1286_.Y
rlabel metal1 2084 3602 2176 3618 0 _1605_.gnd
rlabel metal1 2084 3842 2176 3858 0 _1605_.vdd
rlabel metal2 2093 3693 2107 3707 0 _1605_.A
rlabel metal2 2133 3693 2147 3707 0 _1605_.Y
rlabel metal1 1904 3602 1996 3618 0 _1285_.gnd
rlabel metal1 1904 3842 1996 3858 0 _1285_.vdd
rlabel metal2 1973 3733 1987 3747 0 _1285_.A
rlabel metal2 1933 3733 1947 3747 0 _1285_.B
rlabel metal2 1953 3713 1967 3727 0 _1285_.Y
rlabel metal1 1984 3602 2096 3618 0 _1283_.gnd
rlabel metal1 1984 3842 2096 3858 0 _1283_.vdd
rlabel metal2 1993 3673 2007 3687 0 _1283_.A
rlabel metal2 2013 3693 2027 3707 0 _1283_.B
rlabel metal2 2053 3713 2067 3727 0 _1283_.Y
rlabel metal1 2164 3602 2376 3618 0 CLKBUF1_insert8.gnd
rlabel metal1 2164 3842 2376 3858 0 CLKBUF1_insert8.vdd
rlabel metal2 2333 3713 2347 3727 0 CLKBUF1_insert8.A
rlabel metal2 2193 3713 2207 3727 0 CLKBUF1_insert8.Y
rlabel metal1 2364 3602 2616 3618 0 _1556_.gnd
rlabel metal1 2364 3842 2616 3858 0 _1556_.vdd
rlabel metal2 2453 3693 2467 3707 0 _1556_.D
rlabel metal2 2493 3693 2507 3707 0 _1556_.CLK
rlabel metal2 2573 3693 2587 3707 0 _1556_.Q
rlabel metal1 2604 3602 2716 3618 0 _1275_.gnd
rlabel metal1 2604 3842 2716 3858 0 _1275_.vdd
rlabel metal2 2693 3693 2707 3707 0 _1275_.A
rlabel metal2 2673 3713 2687 3727 0 _1275_.B
rlabel metal2 2633 3713 2647 3727 0 _1275_.C
rlabel metal2 2653 3693 2667 3707 0 _1275_.Y
rlabel metal1 2924 3602 3016 3618 0 _1423_.gnd
rlabel metal1 2924 3842 3016 3858 0 _1423_.vdd
rlabel metal2 2953 3693 2967 3707 0 _1423_.B
rlabel metal2 2993 3693 3007 3707 0 _1423_.A
rlabel metal2 2973 3673 2987 3687 0 _1423_.Y
rlabel metal1 2844 3602 2936 3618 0 _1422_.gnd
rlabel metal1 2844 3842 2936 3858 0 _1422_.vdd
rlabel metal2 2873 3693 2887 3707 0 _1422_.B
rlabel metal2 2913 3693 2927 3707 0 _1422_.A
rlabel metal2 2893 3673 2907 3687 0 _1422_.Y
rlabel metal1 2764 3602 2856 3618 0 _1421_.gnd
rlabel metal1 2764 3842 2856 3858 0 _1421_.vdd
rlabel metal2 2793 3693 2807 3707 0 _1421_.B
rlabel metal2 2833 3693 2847 3707 0 _1421_.A
rlabel metal2 2813 3673 2827 3687 0 _1421_.Y
rlabel metal1 2704 3602 2776 3618 0 _1238_.gnd
rlabel metal1 2704 3842 2776 3858 0 _1238_.vdd
rlabel metal2 2753 3673 2767 3687 0 _1238_.A
rlabel metal2 2733 3713 2747 3727 0 _1238_.Y
rlabel metal1 3124 3602 3236 3618 0 _1429_.gnd
rlabel metal1 3124 3842 3236 3858 0 _1429_.vdd
rlabel metal2 3133 3693 3147 3707 0 _1429_.A
rlabel metal2 3153 3713 3167 3727 0 _1429_.B
rlabel metal2 3193 3713 3207 3727 0 _1429_.C
rlabel metal2 3173 3693 3187 3707 0 _1429_.Y
rlabel metal1 3064 3602 3136 3618 0 _1428_.gnd
rlabel metal1 3064 3842 3136 3858 0 _1428_.vdd
rlabel metal2 3113 3673 3127 3687 0 _1428_.A
rlabel metal2 3093 3713 3107 3727 0 _1428_.Y
rlabel metal1 3004 3602 3076 3618 0 _1424_.gnd
rlabel metal1 3004 3842 3076 3858 0 _1424_.vdd
rlabel metal2 3013 3673 3027 3687 0 _1424_.A
rlabel metal2 3033 3713 3047 3727 0 _1424_.Y
rlabel metal1 3324 3602 3436 3618 0 _1439_.gnd
rlabel metal1 3324 3842 3436 3858 0 _1439_.vdd
rlabel metal2 3333 3713 3347 3727 0 _1439_.A
rlabel metal2 3353 3673 3367 3687 0 _1439_.B
rlabel metal2 3373 3713 3387 3727 0 _1439_.C
rlabel metal2 3393 3693 3407 3707 0 _1439_.Y
rlabel metal1 3224 3602 3336 3618 0 _1420_.gnd
rlabel metal1 3224 3842 3336 3858 0 _1420_.vdd
rlabel metal2 3313 3713 3327 3727 0 _1420_.A
rlabel metal2 3293 3673 3307 3687 0 _1420_.B
rlabel metal2 3273 3713 3287 3727 0 _1420_.C
rlabel metal2 3253 3693 3267 3707 0 _1420_.Y
rlabel metal1 3424 3602 3496 3618 0 _1434_.gnd
rlabel metal1 3424 3842 3496 3858 0 _1434_.vdd
rlabel metal2 3433 3673 3447 3687 0 _1434_.A
rlabel metal2 3453 3713 3467 3727 0 _1434_.Y
rlabel metal1 3684 3602 3796 3618 0 _1427_.gnd
rlabel metal1 3684 3842 3796 3858 0 _1427_.vdd
rlabel metal2 3693 3693 3707 3707 0 _1427_.A
rlabel metal2 3713 3713 3727 3727 0 _1427_.B
rlabel metal2 3753 3713 3767 3727 0 _1427_.C
rlabel metal2 3733 3693 3747 3707 0 _1427_.Y
rlabel metal1 3584 3602 3696 3618 0 _1426_.gnd
rlabel metal1 3584 3842 3696 3858 0 _1426_.vdd
rlabel metal2 3593 3693 3607 3707 0 _1426_.A
rlabel metal2 3613 3713 3627 3727 0 _1426_.B
rlabel metal2 3653 3713 3667 3727 0 _1426_.C
rlabel metal2 3633 3693 3647 3707 0 _1426_.Y
rlabel metal1 3484 3602 3596 3618 0 _1425_.gnd
rlabel metal1 3484 3842 3596 3858 0 _1425_.vdd
rlabel metal2 3493 3693 3507 3707 0 _1425_.A
rlabel metal2 3553 3693 3567 3707 0 _1425_.Y
rlabel metal2 3533 3733 3547 3747 0 _1425_.B
rlabel metal1 3784 3602 4036 3618 0 _1570_.gnd
rlabel metal1 3784 3842 4036 3858 0 _1570_.vdd
rlabel metal2 3873 3693 3887 3707 0 _1570_.D
rlabel metal2 3913 3693 3927 3707 0 _1570_.CLK
rlabel metal2 3993 3693 4007 3707 0 _1570_.Q
rlabel metal1 4024 3602 4116 3618 0 BUFX2_insert5.gnd
rlabel metal1 4024 3842 4116 3858 0 BUFX2_insert5.vdd
rlabel metal2 4033 3693 4047 3707 0 BUFX2_insert5.A
rlabel metal2 4073 3693 4087 3707 0 BUFX2_insert5.Y
rlabel metal1 4184 3602 4296 3618 0 _1500_.gnd
rlabel metal1 4184 3842 4296 3858 0 _1500_.vdd
rlabel metal2 4193 3713 4207 3727 0 _1500_.A
rlabel metal2 4213 3673 4227 3687 0 _1500_.B
rlabel metal2 4233 3713 4247 3727 0 _1500_.C
rlabel metal2 4253 3693 4267 3707 0 _1500_.Y
rlabel metal1 4104 3602 4196 3618 0 _1499_.gnd
rlabel metal1 4104 3842 4196 3858 0 _1499_.vdd
rlabel metal2 4133 3693 4147 3707 0 _1499_.B
rlabel metal2 4173 3693 4187 3707 0 _1499_.A
rlabel metal2 4153 3673 4167 3687 0 _1499_.Y
rlabel metal1 4524 3602 4616 3618 0 _1608_.gnd
rlabel metal1 4524 3842 4616 3858 0 _1608_.vdd
rlabel metal2 4533 3693 4547 3707 0 _1608_.A
rlabel metal2 4573 3693 4587 3707 0 _1608_.Y
rlabel metal1 4284 3602 4536 3618 0 _1583_.gnd
rlabel metal1 4284 3842 4536 3858 0 _1583_.vdd
rlabel metal2 4433 3693 4447 3707 0 _1583_.D
rlabel metal2 4393 3693 4407 3707 0 _1583_.CLK
rlabel metal2 4313 3693 4327 3707 0 _1583_.Q
rlabel nsubstratencontact 4756 3848 4756 3848 0 FILL71250x54150.vdd
rlabel metal1 4744 3602 4776 3618 0 FILL71250x54150.gnd
rlabel nsubstratencontact 4736 3848 4736 3848 0 FILL70950x54150.vdd
rlabel metal1 4724 3602 4756 3618 0 FILL70950x54150.gnd
rlabel metal1 4604 3602 4676 3618 0 _1486_.gnd
rlabel metal1 4604 3842 4676 3858 0 _1486_.vdd
rlabel metal2 4653 3673 4667 3687 0 _1486_.A
rlabel metal2 4633 3713 4647 3727 0 _1486_.Y
rlabel metal1 4664 3602 4736 3618 0 _1483_.gnd
rlabel metal1 4664 3842 4736 3858 0 _1483_.vdd
rlabel metal2 4673 3673 4687 3687 0 _1483_.A
rlabel metal2 4693 3713 4707 3727 0 _1483_.Y
rlabel metal1 244 4082 356 4098 0 _1169_.gnd
rlabel metal1 244 3842 356 3858 0 _1169_.vdd
rlabel metal2 333 3993 347 4007 0 _1169_.A
rlabel metal2 313 3973 327 3987 0 _1169_.B
rlabel metal2 273 3973 287 3987 0 _1169_.C
rlabel metal2 293 3993 307 4007 0 _1169_.Y
rlabel metal1 4 4082 96 4098 0 _1221_.gnd
rlabel metal1 4 3842 96 3858 0 _1221_.vdd
rlabel metal2 73 3953 87 3967 0 _1221_.A
rlabel metal2 33 3953 47 3967 0 _1221_.B
rlabel metal2 53 3973 67 3987 0 _1221_.Y
rlabel metal1 84 4082 176 4098 0 _1172_.gnd
rlabel metal1 84 3842 176 3858 0 _1172_.vdd
rlabel metal2 93 3953 107 3967 0 _1172_.A
rlabel metal2 133 3953 147 3967 0 _1172_.B
rlabel metal2 113 3973 127 3987 0 _1172_.Y
rlabel metal1 164 4082 256 4098 0 _1171_.gnd
rlabel metal1 164 3842 256 3858 0 _1171_.vdd
rlabel metal2 233 3953 247 3967 0 _1171_.A
rlabel metal2 193 3953 207 3967 0 _1171_.B
rlabel metal2 213 3973 227 3987 0 _1171_.Y
rlabel metal1 524 4082 616 4098 0 _1204_.gnd
rlabel metal1 524 3842 616 3858 0 _1204_.vdd
rlabel metal2 533 3953 547 3967 0 _1204_.A
rlabel metal2 573 3953 587 3967 0 _1204_.B
rlabel metal2 553 3973 567 3987 0 _1204_.Y
rlabel metal1 344 4082 456 4098 0 _1222_.gnd
rlabel metal1 344 3842 456 3858 0 _1222_.vdd
rlabel metal2 353 3973 367 3987 0 _1222_.A
rlabel metal2 373 4013 387 4027 0 _1222_.B
rlabel metal2 393 3973 407 3987 0 _1222_.C
rlabel metal2 413 3993 427 4007 0 _1222_.Y
rlabel metal1 444 4082 536 4098 0 _1168_.gnd
rlabel metal1 444 3842 536 3858 0 _1168_.vdd
rlabel metal2 473 3993 487 4007 0 _1168_.B
rlabel metal2 513 3993 527 4007 0 _1168_.A
rlabel metal2 493 4013 507 4027 0 _1168_.Y
rlabel metal1 604 4082 716 4098 0 _1205_.gnd
rlabel metal1 604 3842 716 3858 0 _1205_.vdd
rlabel metal2 613 3993 627 4007 0 _1205_.A
rlabel metal2 633 3973 647 3987 0 _1205_.B
rlabel metal2 673 3973 687 3987 0 _1205_.C
rlabel metal2 653 3993 667 4007 0 _1205_.Y
rlabel metal1 704 4082 816 4098 0 _1220_.gnd
rlabel metal1 704 3842 816 3858 0 _1220_.vdd
rlabel metal2 793 3973 807 3987 0 _1220_.A
rlabel metal2 773 3953 787 3967 0 _1220_.B
rlabel metal2 753 3973 767 3987 0 _1220_.C
rlabel metal2 733 3953 747 3967 0 _1220_.Y
rlabel metal1 1004 4082 1116 4098 0 _1228_.gnd
rlabel metal1 1004 3842 1116 3858 0 _1228_.vdd
rlabel metal2 1013 3993 1027 4007 0 _1228_.A
rlabel metal2 1033 3973 1047 3987 0 _1228_.B
rlabel metal2 1073 3973 1087 3987 0 _1228_.C
rlabel metal2 1053 3993 1067 4007 0 _1228_.Y
rlabel metal1 904 4082 1016 4098 0 _1225_.gnd
rlabel metal1 904 3842 1016 3858 0 _1225_.vdd
rlabel metal2 993 3993 1007 4007 0 _1225_.A
rlabel metal2 973 3973 987 3987 0 _1225_.B
rlabel metal2 933 3973 947 3987 0 _1225_.C
rlabel metal2 953 3993 967 4007 0 _1225_.Y
rlabel metal1 804 4082 916 4098 0 _1227_.gnd
rlabel metal1 804 3842 916 3858 0 _1227_.vdd
rlabel metal2 813 3973 827 3987 0 _1227_.A
rlabel metal2 833 3953 847 3967 0 _1227_.B
rlabel metal2 853 3973 867 3987 0 _1227_.C
rlabel metal2 873 3953 887 3967 0 _1227_.Y
rlabel metal1 1104 4082 1176 4098 0 _1224_.gnd
rlabel metal1 1104 3842 1176 3858 0 _1224_.vdd
rlabel metal2 1153 4013 1167 4027 0 _1224_.A
rlabel metal2 1133 3973 1147 3987 0 _1224_.Y
rlabel metal1 1264 4082 1336 4098 0 _1203_.gnd
rlabel metal1 1264 3842 1336 3858 0 _1203_.vdd
rlabel metal2 1273 4013 1287 4027 0 _1203_.A
rlabel metal2 1293 3973 1307 3987 0 _1203_.Y
rlabel metal1 1164 4082 1276 4098 0 _1232_.gnd
rlabel metal1 1164 3842 1276 3858 0 _1232_.vdd
rlabel metal2 1253 3973 1267 3987 0 _1232_.A
rlabel metal2 1233 3953 1247 3967 0 _1232_.B
rlabel metal2 1213 3973 1227 3987 0 _1232_.C
rlabel metal2 1193 3953 1207 3967 0 _1232_.Y
rlabel metal1 1324 4082 1436 4098 0 _1226_.gnd
rlabel metal1 1324 3842 1436 3858 0 _1226_.vdd
rlabel metal2 1333 3973 1347 3987 0 _1226_.A
rlabel metal2 1353 3953 1367 3967 0 _1226_.B
rlabel metal2 1373 3973 1387 3987 0 _1226_.C
rlabel metal2 1393 3953 1407 3967 0 _1226_.Y
rlabel metal1 1524 4082 1616 4098 0 _1265_.gnd
rlabel metal1 1524 3842 1616 3858 0 _1265_.vdd
rlabel metal2 1533 3953 1547 3967 0 _1265_.A
rlabel metal2 1573 3953 1587 3967 0 _1265_.B
rlabel metal2 1553 3973 1567 3987 0 _1265_.Y
rlabel metal1 1604 4082 1696 4098 0 _1300_.gnd
rlabel metal1 1604 3842 1696 3858 0 _1300_.vdd
rlabel metal2 1633 3993 1647 4007 0 _1300_.B
rlabel metal2 1673 3993 1687 4007 0 _1300_.A
rlabel metal2 1653 4013 1667 4027 0 _1300_.Y
rlabel metal1 1424 4082 1536 4098 0 _1266_.gnd
rlabel metal1 1424 3842 1536 3858 0 _1266_.vdd
rlabel metal2 1433 3973 1447 3987 0 _1266_.A
rlabel metal2 1453 3953 1467 3967 0 _1266_.B
rlabel metal2 1473 3973 1487 3987 0 _1266_.C
rlabel metal2 1493 3953 1507 3967 0 _1266_.Y
rlabel metal1 1784 4082 1896 4098 0 _1301_.gnd
rlabel metal1 1784 3842 1896 3858 0 _1301_.vdd
rlabel metal2 1873 3993 1887 4007 0 _1301_.A
rlabel metal2 1853 3973 1867 3987 0 _1301_.B
rlabel metal2 1813 3973 1827 3987 0 _1301_.C
rlabel metal2 1833 3993 1847 4007 0 _1301_.Y
rlabel metal1 1684 4082 1796 4098 0 _1287_.gnd
rlabel metal1 1684 3842 1796 3858 0 _1287_.vdd
rlabel metal2 1773 3993 1787 4007 0 _1287_.A
rlabel metal2 1713 3993 1727 4007 0 _1287_.Y
rlabel metal2 1733 3953 1747 3967 0 _1287_.B
rlabel metal1 2024 4082 2136 4098 0 _1273_.gnd
rlabel metal1 2024 3842 2136 3858 0 _1273_.vdd
rlabel metal2 2033 3993 2047 4007 0 _1273_.A
rlabel metal2 2053 3973 2067 3987 0 _1273_.B
rlabel metal2 2093 3973 2107 3987 0 _1273_.C
rlabel metal2 2073 3993 2087 4007 0 _1273_.Y
rlabel metal1 1884 4082 1976 4098 0 _1297_.gnd
rlabel metal1 1884 3842 1976 3858 0 _1297_.vdd
rlabel metal2 1933 3993 1947 4007 0 _1297_.B
rlabel metal2 1893 3993 1907 4007 0 _1297_.A
rlabel metal2 1913 4013 1927 4027 0 _1297_.Y
rlabel metal1 1964 4082 2036 4098 0 _1298_.gnd
rlabel metal1 1964 3842 2036 3858 0 _1298_.vdd
rlabel metal2 2013 4013 2027 4027 0 _1298_.A
rlabel metal2 1993 3973 2007 3987 0 _1298_.Y
rlabel metal1 2124 4082 2196 4098 0 _1272_.gnd
rlabel metal1 2124 3842 2196 3858 0 _1272_.vdd
rlabel metal2 2133 4013 2147 4027 0 _1272_.A
rlabel metal2 2153 3973 2167 3987 0 _1272_.Y
rlabel metal1 2364 4082 2456 4098 0 _1603_.gnd
rlabel metal1 2364 3842 2456 3858 0 _1603_.vdd
rlabel metal2 2373 3993 2387 4007 0 _1603_.A
rlabel metal2 2413 3993 2427 4007 0 _1603_.Y
rlabel metal1 2184 4082 2276 4098 0 _1268_.gnd
rlabel metal1 2184 3842 2276 3858 0 _1268_.vdd
rlabel metal2 2193 3953 2207 3967 0 _1268_.A
rlabel metal2 2233 3953 2247 3967 0 _1268_.B
rlabel metal2 2213 3973 2227 3987 0 _1268_.Y
rlabel metal1 2264 4082 2376 4098 0 _1274_.gnd
rlabel metal1 2264 3842 2376 3858 0 _1274_.vdd
rlabel metal2 2273 3973 2287 3987 0 _1274_.A
rlabel metal2 2293 3953 2307 3967 0 _1274_.B
rlabel metal2 2313 3973 2327 3987 0 _1274_.C
rlabel metal2 2333 3953 2347 3967 0 _1274_.Y
rlabel metal1 2444 4082 2656 4098 0 CLKBUF1_insert12.gnd
rlabel metal1 2444 3842 2656 3858 0 CLKBUF1_insert12.vdd
rlabel metal2 2473 3973 2487 3987 0 CLKBUF1_insert12.A
rlabel metal2 2613 3973 2627 3987 0 CLKBUF1_insert12.Y
rlabel metal1 2644 4082 2896 4098 0 _1540_.gnd
rlabel metal1 2644 3842 2896 3858 0 _1540_.vdd
rlabel metal2 2733 3993 2747 4007 0 _1540_.D
rlabel metal2 2773 3993 2787 4007 0 _1540_.CLK
rlabel metal2 2853 3993 2867 4007 0 _1540_.Q
rlabel metal1 2884 4082 2956 4098 0 _833_.gnd
rlabel metal1 2884 3842 2956 3858 0 _833_.vdd
rlabel metal2 2893 4013 2907 4027 0 _833_.A
rlabel metal2 2913 3973 2927 3987 0 _833_.Y
rlabel metal1 2944 4082 3056 4098 0 _835_.gnd
rlabel metal1 2944 3842 3056 3858 0 _835_.vdd
rlabel metal2 2953 3993 2967 4007 0 _835_.A
rlabel metal2 2973 3973 2987 3987 0 _835_.B
rlabel metal2 3013 3973 3027 3987 0 _835_.C
rlabel metal2 2993 3993 3007 4007 0 _835_.Y
rlabel metal1 3124 4082 3216 4098 0 _834_.gnd
rlabel metal1 3124 3842 3216 3858 0 _834_.vdd
rlabel metal2 3133 3953 3147 3967 0 _834_.A
rlabel metal2 3173 3953 3187 3967 0 _834_.B
rlabel metal2 3153 3973 3167 3987 0 _834_.Y
rlabel metal1 3204 4082 3316 4098 0 _1408_.gnd
rlabel metal1 3204 3842 3316 3858 0 _1408_.vdd
rlabel metal2 3293 3973 3307 3987 0 _1408_.A
rlabel metal2 3273 4013 3287 4027 0 _1408_.B
rlabel metal2 3253 3973 3267 3987 0 _1408_.C
rlabel metal2 3233 3993 3247 4007 0 _1408_.Y
rlabel metal1 3044 4082 3136 4098 0 _1403_.gnd
rlabel metal1 3044 3842 3136 3858 0 _1403_.vdd
rlabel metal2 3093 3993 3107 4007 0 _1403_.B
rlabel metal2 3053 3993 3067 4007 0 _1403_.A
rlabel metal2 3073 4013 3087 4027 0 _1403_.Y
rlabel metal1 3404 4082 3496 4098 0 _1433_.gnd
rlabel metal1 3404 3842 3496 3858 0 _1433_.vdd
rlabel metal2 3433 3993 3447 4007 0 _1433_.B
rlabel metal2 3473 3993 3487 4007 0 _1433_.A
rlabel metal2 3453 4013 3467 4027 0 _1433_.Y
rlabel metal1 3304 4082 3416 4098 0 _1417_.gnd
rlabel metal1 3304 3842 3416 3858 0 _1417_.vdd
rlabel metal2 3313 3993 3327 4007 0 _1417_.A
rlabel metal2 3373 3993 3387 4007 0 _1417_.Y
rlabel metal2 3353 3953 3367 3967 0 _1417_.B
rlabel metal1 3544 4082 3796 4098 0 _1582_.gnd
rlabel metal1 3544 3842 3796 3858 0 _1582_.vdd
rlabel metal2 3693 3993 3707 4007 0 _1582_.D
rlabel metal2 3653 3993 3667 4007 0 _1582_.CLK
rlabel metal2 3573 3993 3587 4007 0 _1582_.Q
rlabel metal1 3484 4082 3556 4098 0 _1432_.gnd
rlabel metal1 3484 3842 3556 3858 0 _1432_.vdd
rlabel metal2 3533 4013 3547 4027 0 _1432_.A
rlabel metal2 3513 3973 3527 3987 0 _1432_.Y
rlabel metal1 3784 4082 3896 4098 0 _1498_.gnd
rlabel metal1 3784 3842 3896 3858 0 _1498_.vdd
rlabel metal2 3873 3973 3887 3987 0 _1498_.A
rlabel metal2 3853 4013 3867 4027 0 _1498_.B
rlabel metal2 3833 3973 3847 3987 0 _1498_.C
rlabel metal2 3813 3993 3827 4007 0 _1498_.Y
rlabel metal1 3884 4082 3976 4098 0 _1497_.gnd
rlabel metal1 3884 3842 3976 3858 0 _1497_.vdd
rlabel metal2 3933 3993 3947 4007 0 _1497_.B
rlabel metal2 3893 3993 3907 4007 0 _1497_.A
rlabel metal2 3913 4013 3927 4027 0 _1497_.Y
rlabel metal1 3964 4082 4056 4098 0 _1413_.gnd
rlabel metal1 3964 3842 4056 3858 0 _1413_.vdd
rlabel metal2 3993 3993 4007 4007 0 _1413_.B
rlabel metal2 4033 3993 4047 4007 0 _1413_.A
rlabel metal2 4013 4013 4027 4027 0 _1413_.Y
rlabel metal1 4244 4082 4356 4098 0 _1415_.gnd
rlabel metal1 4244 3842 4356 3858 0 _1415_.vdd
rlabel metal2 4333 3993 4347 4007 0 _1415_.A
rlabel metal2 4313 3973 4327 3987 0 _1415_.B
rlabel metal2 4273 3973 4287 3987 0 _1415_.C
rlabel metal2 4293 3993 4307 4007 0 _1415_.Y
rlabel metal1 4144 4082 4256 4098 0 _1414_.gnd
rlabel metal1 4144 3842 4256 3858 0 _1414_.vdd
rlabel metal2 4153 3993 4167 4007 0 _1414_.A
rlabel metal2 4173 3973 4187 3987 0 _1414_.B
rlabel metal2 4213 3973 4227 3987 0 _1414_.C
rlabel metal2 4193 3993 4207 4007 0 _1414_.Y
rlabel metal1 4044 4082 4156 4098 0 _1412_.gnd
rlabel metal1 4044 3842 4156 3858 0 _1412_.vdd
rlabel metal2 4053 3993 4067 4007 0 _1412_.A
rlabel metal2 4113 3993 4127 4007 0 _1412_.Y
rlabel metal2 4093 3953 4107 3967 0 _1412_.B
rlabel metal1 4404 4082 4656 4098 0 _1569_.gnd
rlabel metal1 4404 3842 4656 3858 0 _1569_.vdd
rlabel metal2 4553 3993 4567 4007 0 _1569_.D
rlabel metal2 4513 3993 4527 4007 0 _1569_.CLK
rlabel metal2 4433 3993 4447 4007 0 _1569_.Q
rlabel metal1 4344 4082 4416 4098 0 _769_.gnd
rlabel metal1 4344 3842 4416 3858 0 _769_.vdd
rlabel metal2 4393 4013 4407 4027 0 _769_.A
rlabel metal2 4373 3973 4387 3987 0 _769_.Y
rlabel nsubstratencontact 4764 3852 4764 3852 0 FILL71250x57750.vdd
rlabel metal1 4744 4082 4776 4098 0 FILL71250x57750.gnd
rlabel nsubstratencontact 4744 3852 4744 3852 0 FILL70950x57750.vdd
rlabel metal1 4724 4082 4756 4098 0 FILL70950x57750.gnd
rlabel nsubstratencontact 4724 3852 4724 3852 0 FILL70650x57750.vdd
rlabel metal1 4704 4082 4736 4098 0 FILL70650x57750.gnd
rlabel metal1 4644 4082 4716 4098 0 _1479_.gnd
rlabel metal1 4644 3842 4716 3858 0 _1479_.vdd
rlabel metal2 4653 4013 4667 4027 0 _1479_.A
rlabel metal2 4673 3973 4687 3987 0 _1479_.Y
rlabel metal1 184 4082 276 4098 0 _1174_.gnd
rlabel metal1 184 4322 276 4338 0 _1174_.vdd
rlabel metal2 253 4213 267 4227 0 _1174_.A
rlabel metal2 213 4213 227 4227 0 _1174_.B
rlabel metal2 233 4193 247 4207 0 _1174_.Y
rlabel metal1 4 4082 96 4098 0 _1173_.gnd
rlabel metal1 4 4322 96 4338 0 _1173_.vdd
rlabel metal2 73 4213 87 4227 0 _1173_.A
rlabel metal2 33 4213 47 4227 0 _1173_.B
rlabel metal2 53 4193 67 4207 0 _1173_.Y
rlabel metal1 84 4082 196 4098 0 _1179_.gnd
rlabel metal1 84 4322 196 4338 0 _1179_.vdd
rlabel metal2 93 4193 107 4207 0 _1179_.A
rlabel metal2 113 4153 127 4167 0 _1179_.B
rlabel metal2 133 4193 147 4207 0 _1179_.C
rlabel metal2 153 4173 167 4187 0 _1179_.Y
rlabel metal1 264 4082 356 4098 0 _1178_.gnd
rlabel metal1 264 4322 356 4338 0 _1178_.vdd
rlabel metal2 293 4173 307 4187 0 _1178_.B
rlabel metal2 333 4173 347 4187 0 _1178_.A
rlabel metal2 313 4153 327 4167 0 _1178_.Y
rlabel metal1 444 4082 556 4098 0 _1183_.gnd
rlabel metal1 444 4322 556 4338 0 _1183_.vdd
rlabel metal2 453 4173 467 4187 0 _1183_.A
rlabel metal2 473 4193 487 4207 0 _1183_.B
rlabel metal2 513 4193 527 4207 0 _1183_.C
rlabel metal2 493 4173 507 4187 0 _1183_.Y
rlabel metal1 344 4082 456 4098 0 _1180_.gnd
rlabel metal1 344 4322 456 4338 0 _1180_.vdd
rlabel metal2 433 4173 447 4187 0 _1180_.A
rlabel metal2 413 4193 427 4207 0 _1180_.B
rlabel metal2 373 4193 387 4207 0 _1180_.C
rlabel metal2 393 4173 407 4187 0 _1180_.Y
rlabel metal1 604 4082 716 4098 0 _1187_.gnd
rlabel metal1 604 4322 716 4338 0 _1187_.vdd
rlabel metal2 693 4193 707 4207 0 _1187_.A
rlabel metal2 673 4153 687 4167 0 _1187_.B
rlabel metal2 653 4193 667 4207 0 _1187_.C
rlabel metal2 633 4173 647 4187 0 _1187_.Y
rlabel metal1 704 4082 776 4098 0 _1186_.gnd
rlabel metal1 704 4322 776 4338 0 _1186_.vdd
rlabel metal2 753 4153 767 4167 0 _1186_.A
rlabel metal2 733 4193 747 4207 0 _1186_.Y
rlabel metal1 544 4082 616 4098 0 _1143_.gnd
rlabel metal1 544 4322 616 4338 0 _1143_.vdd
rlabel metal2 593 4153 607 4167 0 _1143_.A
rlabel metal2 573 4193 587 4207 0 _1143_.Y
rlabel metal1 764 4082 876 4098 0 _1184_.gnd
rlabel metal1 764 4322 876 4338 0 _1184_.vdd
rlabel metal2 773 4193 787 4207 0 _1184_.A
rlabel metal2 793 4213 807 4227 0 _1184_.B
rlabel metal2 813 4193 827 4207 0 _1184_.C
rlabel metal2 833 4213 847 4227 0 _1184_.Y
rlabel metal1 984 4082 1096 4098 0 _1231_.gnd
rlabel metal1 984 4322 1096 4338 0 _1231_.vdd
rlabel metal2 1073 4193 1087 4207 0 _1231_.A
rlabel metal2 1053 4213 1067 4227 0 _1231_.B
rlabel metal2 1033 4193 1047 4207 0 _1231_.C
rlabel metal2 1013 4213 1027 4227 0 _1231_.Y
rlabel metal1 864 4082 996 4098 0 _1233_.gnd
rlabel metal1 864 4322 996 4338 0 _1233_.vdd
rlabel metal2 973 4173 987 4187 0 _1233_.A
rlabel metal2 953 4193 967 4207 0 _1233_.B
rlabel metal2 893 4173 907 4187 0 _1233_.C
rlabel metal2 913 4193 927 4207 0 _1233_.D
rlabel metal2 933 4173 947 4187 0 _1233_.Y
rlabel metal1 1184 4082 1276 4098 0 _1246_.gnd
rlabel metal1 1184 4322 1276 4338 0 _1246_.vdd
rlabel metal2 1253 4213 1267 4227 0 _1246_.A
rlabel metal2 1213 4213 1227 4227 0 _1246_.B
rlabel metal2 1233 4193 1247 4207 0 _1246_.Y
rlabel metal1 1264 4082 1376 4098 0 _1264_.gnd
rlabel metal1 1264 4322 1376 4338 0 _1264_.vdd
rlabel metal2 1353 4193 1367 4207 0 _1264_.A
rlabel metal2 1333 4213 1347 4227 0 _1264_.B
rlabel metal2 1313 4193 1327 4207 0 _1264_.C
rlabel metal2 1293 4213 1307 4227 0 _1264_.Y
rlabel metal1 1084 4082 1196 4098 0 _1229_.gnd
rlabel metal1 1084 4322 1196 4338 0 _1229_.vdd
rlabel metal2 1093 4193 1107 4207 0 _1229_.A
rlabel metal2 1113 4213 1127 4227 0 _1229_.B
rlabel metal2 1133 4193 1147 4207 0 _1229_.C
rlabel metal2 1153 4213 1167 4227 0 _1229_.Y
rlabel metal1 1364 4082 1456 4098 0 _1267_.gnd
rlabel metal1 1364 4322 1456 4338 0 _1267_.vdd
rlabel metal2 1433 4213 1447 4227 0 _1267_.A
rlabel metal2 1393 4213 1407 4227 0 _1267_.B
rlabel metal2 1413 4193 1427 4207 0 _1267_.Y
rlabel metal1 1544 4082 1636 4098 0 _1299_.gnd
rlabel metal1 1544 4322 1636 4338 0 _1299_.vdd
rlabel metal2 1573 4173 1587 4187 0 _1299_.B
rlabel metal2 1613 4173 1627 4187 0 _1299_.A
rlabel metal2 1593 4153 1607 4167 0 _1299_.Y
rlabel metal1 1444 4082 1556 4098 0 _1296_.gnd
rlabel metal1 1444 4322 1556 4338 0 _1296_.vdd
rlabel metal2 1453 4193 1467 4207 0 _1296_.A
rlabel metal2 1473 4213 1487 4227 0 _1296_.B
rlabel metal2 1493 4193 1507 4207 0 _1296_.C
rlabel metal2 1513 4213 1527 4227 0 _1296_.Y
rlabel metal1 1704 4082 1816 4098 0 _1291_.gnd
rlabel metal1 1704 4322 1816 4338 0 _1291_.vdd
rlabel metal2 1713 4173 1727 4187 0 _1291_.A
rlabel metal2 1733 4193 1747 4207 0 _1291_.B
rlabel metal2 1773 4193 1787 4207 0 _1291_.C
rlabel metal2 1753 4173 1767 4187 0 _1291_.Y
rlabel metal1 1804 4082 1896 4098 0 _1292_.gnd
rlabel metal1 1804 4322 1896 4338 0 _1292_.vdd
rlabel metal2 1873 4213 1887 4227 0 _1292_.A
rlabel metal2 1833 4213 1847 4227 0 _1292_.B
rlabel metal2 1853 4193 1867 4207 0 _1292_.Y
rlabel metal1 1624 4082 1716 4098 0 _1288_.gnd
rlabel metal1 1624 4322 1716 4338 0 _1288_.vdd
rlabel metal2 1653 4173 1667 4187 0 _1288_.B
rlabel metal2 1693 4173 1707 4187 0 _1288_.A
rlabel metal2 1673 4153 1687 4167 0 _1288_.Y
rlabel metal1 1884 4082 1956 4098 0 _1289_.gnd
rlabel metal1 1884 4322 1956 4338 0 _1289_.vdd
rlabel metal2 1893 4153 1907 4167 0 _1289_.A
rlabel metal2 1913 4193 1927 4207 0 _1289_.Y
rlabel metal1 2044 4082 2156 4098 0 _1293_.gnd
rlabel metal1 2044 4322 2156 4338 0 _1293_.vdd
rlabel metal2 2053 4193 2067 4207 0 _1293_.A
rlabel metal2 2073 4213 2087 4227 0 _1293_.B
rlabel metal2 2093 4193 2107 4207 0 _1293_.C
rlabel metal2 2113 4213 2127 4227 0 _1293_.Y
rlabel metal1 1944 4082 2056 4098 0 _1290_.gnd
rlabel metal1 1944 4322 2056 4338 0 _1290_.vdd
rlabel metal2 1953 4193 1967 4207 0 _1290_.A
rlabel metal2 1973 4213 1987 4227 0 _1290_.B
rlabel metal2 1993 4193 2007 4207 0 _1290_.C
rlabel metal2 2013 4213 2027 4227 0 _1290_.Y
rlabel metal1 2384 4082 2476 4098 0 _1604_.gnd
rlabel metal1 2384 4322 2476 4338 0 _1604_.vdd
rlabel metal2 2393 4173 2407 4187 0 _1604_.A
rlabel metal2 2433 4173 2447 4187 0 _1604_.Y
rlabel metal1 2144 4082 2396 4098 0 _1554_.gnd
rlabel metal1 2144 4322 2396 4338 0 _1554_.vdd
rlabel metal2 2233 4173 2247 4187 0 _1554_.D
rlabel metal2 2273 4173 2287 4187 0 _1554_.CLK
rlabel metal2 2353 4173 2367 4187 0 _1554_.Q
rlabel metal1 2604 4082 2856 4098 0 _1538_.gnd
rlabel metal1 2604 4322 2856 4338 0 _1538_.vdd
rlabel metal2 2753 4173 2767 4187 0 _1538_.D
rlabel metal2 2713 4173 2727 4187 0 _1538_.CLK
rlabel metal2 2633 4173 2647 4187 0 _1538_.Q
rlabel metal1 2524 4082 2616 4098 0 _1401_.gnd
rlabel metal1 2524 4322 2616 4338 0 _1401_.vdd
rlabel metal2 2553 4173 2567 4187 0 _1401_.B
rlabel metal2 2593 4173 2607 4187 0 _1401_.A
rlabel metal2 2573 4153 2587 4167 0 _1401_.Y
rlabel metal1 2464 4082 2536 4098 0 _1136_.gnd
rlabel metal1 2464 4322 2536 4338 0 _1136_.vdd
rlabel metal2 2513 4153 2527 4167 0 _1136_.A
rlabel metal2 2493 4193 2507 4207 0 _1136_.Y
rlabel metal1 2904 4082 2996 4098 0 _1402_.gnd
rlabel metal1 2904 4322 2996 4338 0 _1402_.vdd
rlabel metal2 2933 4173 2947 4187 0 _1402_.B
rlabel metal2 2973 4173 2987 4187 0 _1402_.A
rlabel metal2 2953 4153 2967 4167 0 _1402_.Y
rlabel metal1 2844 4082 2916 4098 0 _827_.gnd
rlabel metal1 2844 4322 2916 4338 0 _827_.vdd
rlabel metal2 2853 4153 2867 4167 0 _827_.A
rlabel metal2 2873 4193 2887 4207 0 _827_.Y
rlabel metal1 2984 4082 3096 4098 0 _829_.gnd
rlabel metal1 2984 4322 3096 4338 0 _829_.vdd
rlabel metal2 2993 4173 3007 4187 0 _829_.A
rlabel metal2 3013 4193 3027 4207 0 _829_.B
rlabel metal2 3053 4193 3067 4207 0 _829_.C
rlabel metal2 3033 4173 3047 4187 0 _829_.Y
rlabel metal1 3164 4082 3256 4098 0 _1294_.gnd
rlabel metal1 3164 4322 3256 4338 0 _1294_.vdd
rlabel metal2 3233 4213 3247 4227 0 _1294_.A
rlabel metal2 3193 4213 3207 4227 0 _1294_.B
rlabel metal2 3213 4193 3227 4207 0 _1294_.Y
rlabel metal1 3084 4082 3176 4098 0 _828_.gnd
rlabel metal1 3084 4322 3176 4338 0 _828_.vdd
rlabel metal2 3093 4213 3107 4227 0 _828_.A
rlabel metal2 3133 4213 3147 4227 0 _828_.B
rlabel metal2 3113 4193 3127 4207 0 _828_.Y
rlabel metal1 3404 4082 3656 4098 0 _1557_.gnd
rlabel metal1 3404 4322 3656 4338 0 _1557_.vdd
rlabel metal2 3493 4173 3507 4187 0 _1557_.D
rlabel metal2 3533 4173 3547 4187 0 _1557_.CLK
rlabel metal2 3613 4173 3627 4187 0 _1557_.Q
rlabel metal1 3244 4082 3336 4098 0 _1276_.gnd
rlabel metal1 3244 4322 3336 4338 0 _1276_.vdd
rlabel metal2 3313 4213 3327 4227 0 _1276_.A
rlabel metal2 3273 4213 3287 4227 0 _1276_.B
rlabel metal2 3293 4193 3307 4207 0 _1276_.Y
rlabel metal1 3324 4082 3416 4098 0 _1411_.gnd
rlabel metal1 3324 4322 3416 4338 0 _1411_.vdd
rlabel metal2 3373 4173 3387 4187 0 _1411_.B
rlabel metal2 3333 4173 3347 4187 0 _1411_.A
rlabel metal2 3353 4153 3367 4167 0 _1411_.Y
rlabel metal1 3644 4082 3736 4098 0 _1431_.gnd
rlabel metal1 3644 4322 3736 4338 0 _1431_.vdd
rlabel metal2 3713 4213 3727 4227 0 _1431_.A
rlabel metal2 3673 4213 3687 4227 0 _1431_.B
rlabel metal2 3693 4193 3707 4207 0 _1431_.Y
rlabel metal1 3724 4082 3816 4098 0 _1430_.gnd
rlabel metal1 3724 4322 3816 4338 0 _1430_.vdd
rlabel metal2 3773 4173 3787 4187 0 _1430_.B
rlabel metal2 3733 4173 3747 4187 0 _1430_.A
rlabel metal2 3753 4153 3767 4167 0 _1430_.Y
rlabel metal1 3804 4082 4056 4098 0 _1581_.gnd
rlabel metal1 3804 4322 4056 4338 0 _1581_.vdd
rlabel metal2 3953 4173 3967 4187 0 _1581_.D
rlabel metal2 3913 4173 3927 4187 0 _1581_.CLK
rlabel metal2 3833 4173 3847 4187 0 _1581_.Q
rlabel metal1 4224 4082 4316 4098 0 _1607_.gnd
rlabel metal1 4224 4322 4316 4338 0 _1607_.vdd
rlabel metal2 4233 4173 4247 4187 0 _1607_.A
rlabel metal2 4273 4173 4287 4187 0 _1607_.Y
rlabel metal1 4124 4082 4236 4098 0 _1496_.gnd
rlabel metal1 4124 4322 4236 4338 0 _1496_.vdd
rlabel metal2 4213 4193 4227 4207 0 _1496_.A
rlabel metal2 4193 4153 4207 4167 0 _1496_.B
rlabel metal2 4173 4193 4187 4207 0 _1496_.C
rlabel metal2 4153 4173 4167 4187 0 _1496_.Y
rlabel metal1 4044 4082 4136 4098 0 _1495_.gnd
rlabel metal1 4044 4322 4136 4338 0 _1495_.vdd
rlabel metal2 4093 4173 4107 4187 0 _1495_.B
rlabel metal2 4053 4173 4067 4187 0 _1495_.A
rlabel metal2 4073 4153 4087 4167 0 _1495_.Y
rlabel metal1 4484 4082 4736 4098 0 _1580_.gnd
rlabel metal1 4484 4322 4736 4338 0 _1580_.vdd
rlabel metal2 4633 4173 4647 4187 0 _1580_.D
rlabel metal2 4593 4173 4607 4187 0 _1580_.CLK
rlabel metal2 4513 4173 4527 4187 0 _1580_.Q
rlabel metal1 4384 4082 4496 4098 0 _1494_.gnd
rlabel metal1 4384 4322 4496 4338 0 _1494_.vdd
rlabel metal2 4473 4193 4487 4207 0 _1494_.A
rlabel metal2 4453 4153 4467 4167 0 _1494_.B
rlabel metal2 4433 4193 4447 4207 0 _1494_.C
rlabel metal2 4413 4173 4427 4187 0 _1494_.Y
rlabel metal1 4304 4082 4396 4098 0 _1493_.gnd
rlabel metal1 4304 4322 4396 4338 0 _1493_.vdd
rlabel metal2 4333 4173 4347 4187 0 _1493_.B
rlabel metal2 4373 4173 4387 4187 0 _1493_.A
rlabel metal2 4353 4153 4367 4167 0 _1493_.Y
rlabel nsubstratencontact 4756 4328 4756 4328 0 FILL71250x61350.vdd
rlabel metal1 4744 4082 4776 4098 0 FILL71250x61350.gnd
rlabel nsubstratencontact 4736 4328 4736 4328 0 FILL70950x61350.vdd
rlabel metal1 4724 4082 4756 4098 0 FILL70950x61350.gnd
rlabel metal1 4 4562 116 4578 0 _1200_.gnd
rlabel metal1 4 4322 116 4338 0 _1200_.vdd
rlabel metal2 93 4453 107 4467 0 _1200_.A
rlabel metal2 73 4493 87 4507 0 _1200_.B
rlabel metal2 53 4453 67 4467 0 _1200_.C
rlabel metal2 33 4473 47 4487 0 _1200_.Y
rlabel metal1 104 4562 216 4578 0 _1182_.gnd
rlabel metal1 104 4322 216 4338 0 _1182_.vdd
rlabel metal2 193 4453 207 4467 0 _1182_.A
rlabel metal2 173 4433 187 4447 0 _1182_.B
rlabel metal2 153 4453 167 4467 0 _1182_.C
rlabel metal2 133 4433 147 4447 0 _1182_.Y
rlabel metal1 204 4562 316 4578 0 _1175_.gnd
rlabel metal1 204 4322 316 4338 0 _1175_.vdd
rlabel metal2 213 4453 227 4467 0 _1175_.A
rlabel metal2 233 4433 247 4447 0 _1175_.B
rlabel metal2 253 4453 267 4467 0 _1175_.C
rlabel metal2 273 4433 287 4447 0 _1175_.Y
rlabel metal1 504 4562 616 4578 0 _1201_.gnd
rlabel metal1 504 4322 616 4338 0 _1201_.vdd
rlabel metal2 513 4473 527 4487 0 _1201_.A
rlabel metal2 533 4453 547 4467 0 _1201_.B
rlabel metal2 573 4453 587 4467 0 _1201_.C
rlabel metal2 553 4473 567 4487 0 _1201_.Y
rlabel metal1 404 4562 516 4578 0 _1188_.gnd
rlabel metal1 404 4322 516 4338 0 _1188_.vdd
rlabel metal2 413 4453 427 4467 0 _1188_.A
rlabel metal2 433 4493 447 4507 0 _1188_.B
rlabel metal2 453 4453 467 4467 0 _1188_.C
rlabel metal2 473 4473 487 4487 0 _1188_.Y
rlabel metal1 304 4562 416 4578 0 _1181_.gnd
rlabel metal1 304 4322 416 4338 0 _1181_.vdd
rlabel metal2 393 4453 407 4467 0 _1181_.A
rlabel metal2 373 4433 387 4447 0 _1181_.B
rlabel metal2 353 4453 367 4467 0 _1181_.C
rlabel metal2 333 4433 347 4447 0 _1181_.Y
rlabel metal1 604 4562 716 4578 0 _1189_.gnd
rlabel metal1 604 4322 716 4338 0 _1189_.vdd
rlabel metal2 613 4473 627 4487 0 _1189_.A
rlabel metal2 633 4453 647 4467 0 _1189_.B
rlabel metal2 673 4453 687 4467 0 _1189_.C
rlabel metal2 653 4473 667 4487 0 _1189_.Y
rlabel metal1 704 4562 816 4578 0 _1185_.gnd
rlabel metal1 704 4322 816 4338 0 _1185_.vdd
rlabel metal2 793 4453 807 4467 0 _1185_.A
rlabel metal2 773 4433 787 4447 0 _1185_.B
rlabel metal2 753 4453 767 4467 0 _1185_.C
rlabel metal2 733 4433 747 4447 0 _1185_.Y
rlabel metal1 904 4562 996 4578 0 _1239_.gnd
rlabel metal1 904 4322 996 4338 0 _1239_.vdd
rlabel metal2 913 4433 927 4447 0 _1239_.A
rlabel metal2 953 4433 967 4447 0 _1239_.B
rlabel metal2 933 4453 947 4467 0 _1239_.Y
rlabel metal1 984 4562 1096 4578 0 _1241_.gnd
rlabel metal1 984 4322 1096 4338 0 _1241_.vdd
rlabel metal2 993 4453 1007 4467 0 _1241_.A
rlabel metal2 1013 4433 1027 4447 0 _1241_.B
rlabel metal2 1033 4453 1047 4467 0 _1241_.C
rlabel metal2 1053 4433 1067 4447 0 _1241_.Y
rlabel metal1 804 4562 916 4578 0 _1240_.gnd
rlabel metal1 804 4322 916 4338 0 _1240_.vdd
rlabel metal2 813 4453 827 4467 0 _1240_.A
rlabel metal2 833 4433 847 4447 0 _1240_.B
rlabel metal2 853 4453 867 4467 0 _1240_.C
rlabel metal2 873 4433 887 4447 0 _1240_.Y
rlabel metal1 1184 4562 1276 4578 0 _1242_.gnd
rlabel metal1 1184 4322 1276 4338 0 _1242_.vdd
rlabel metal2 1253 4433 1267 4447 0 _1242_.A
rlabel metal2 1213 4433 1227 4447 0 _1242_.B
rlabel metal2 1233 4453 1247 4467 0 _1242_.Y
rlabel metal1 1084 4562 1196 4578 0 _1230_.gnd
rlabel metal1 1084 4322 1196 4338 0 _1230_.vdd
rlabel metal2 1093 4453 1107 4467 0 _1230_.A
rlabel metal2 1113 4493 1127 4507 0 _1230_.B
rlabel metal2 1133 4453 1147 4467 0 _1230_.C
rlabel metal2 1153 4473 1167 4487 0 _1230_.Y
rlabel metal1 1264 4562 1356 4578 0 _1234_.gnd
rlabel metal1 1264 4322 1356 4338 0 _1234_.vdd
rlabel metal2 1293 4473 1307 4487 0 _1234_.B
rlabel metal2 1333 4473 1347 4487 0 _1234_.A
rlabel metal2 1313 4493 1327 4507 0 _1234_.Y
rlabel metal1 1344 4562 1456 4578 0 _1244_.gnd
rlabel metal1 1344 4322 1456 4338 0 _1244_.vdd
rlabel metal2 1433 4473 1447 4487 0 _1244_.A
rlabel metal2 1413 4453 1427 4467 0 _1244_.B
rlabel metal2 1373 4453 1387 4467 0 _1244_.C
rlabel metal2 1393 4473 1407 4487 0 _1244_.Y
rlabel metal1 1444 4562 1536 4578 0 _1190_.gnd
rlabel metal1 1444 4322 1536 4338 0 _1190_.vdd
rlabel metal2 1513 4433 1527 4447 0 _1190_.A
rlabel metal2 1473 4433 1487 4447 0 _1190_.B
rlabel metal2 1493 4453 1507 4467 0 _1190_.Y
rlabel metal1 1524 4562 1616 4578 0 _1243_.gnd
rlabel metal1 1524 4322 1616 4338 0 _1243_.vdd
rlabel metal2 1573 4473 1587 4487 0 _1243_.B
rlabel metal2 1533 4473 1547 4487 0 _1243_.A
rlabel metal2 1553 4493 1567 4507 0 _1243_.Y
rlabel metal1 1604 4562 1716 4578 0 _1270_.gnd
rlabel metal1 1604 4322 1716 4338 0 _1270_.vdd
rlabel metal2 1613 4453 1627 4467 0 _1270_.A
rlabel metal2 1633 4433 1647 4447 0 _1270_.B
rlabel metal2 1653 4453 1667 4467 0 _1270_.C
rlabel metal2 1673 4433 1687 4447 0 _1270_.Y
rlabel metal1 1704 4562 1816 4578 0 _1245_.gnd
rlabel metal1 1704 4322 1816 4338 0 _1245_.vdd
rlabel metal2 1793 4453 1807 4467 0 _1245_.A
rlabel metal2 1773 4493 1787 4507 0 _1245_.B
rlabel metal2 1753 4453 1767 4467 0 _1245_.C
rlabel metal2 1733 4473 1747 4487 0 _1245_.Y
rlabel metal1 1804 4562 1876 4578 0 _1198_.gnd
rlabel metal1 1804 4322 1876 4338 0 _1198_.vdd
rlabel metal2 1813 4493 1827 4507 0 _1198_.A
rlabel metal2 1833 4453 1847 4467 0 _1198_.Y
rlabel metal1 1864 4562 1936 4578 0 _1191_.gnd
rlabel metal1 1864 4322 1936 4338 0 _1191_.vdd
rlabel metal2 1913 4493 1927 4507 0 _1191_.A
rlabel metal2 1893 4453 1907 4467 0 _1191_.Y
rlabel metal1 1924 4562 2036 4578 0 _1199_.gnd
rlabel metal1 1924 4322 2036 4338 0 _1199_.vdd
rlabel metal2 1933 4453 1947 4467 0 _1199_.A
rlabel metal2 1953 4493 1967 4507 0 _1199_.B
rlabel metal2 1973 4453 1987 4467 0 _1199_.C
rlabel metal2 1993 4473 2007 4487 0 _1199_.Y
rlabel metal1 2024 4562 2116 4578 0 _1192_.gnd
rlabel metal1 2024 4322 2116 4338 0 _1192_.vdd
rlabel metal2 2073 4473 2087 4487 0 _1192_.B
rlabel metal2 2033 4473 2047 4487 0 _1192_.A
rlabel metal2 2053 4493 2067 4507 0 _1192_.Y
rlabel metal1 2104 4562 2176 4578 0 _1193_.gnd
rlabel metal1 2104 4322 2176 4338 0 _1193_.vdd
rlabel metal2 2113 4493 2127 4507 0 _1193_.A
rlabel metal2 2133 4453 2147 4467 0 _1193_.Y
rlabel metal1 2164 4562 2276 4578 0 _1194_.gnd
rlabel metal1 2164 4322 2276 4338 0 _1194_.vdd
rlabel metal2 2173 4473 2187 4487 0 _1194_.A
rlabel metal2 2193 4453 2207 4467 0 _1194_.B
rlabel metal2 2233 4453 2247 4467 0 _1194_.C
rlabel metal2 2213 4473 2227 4487 0 _1194_.Y
rlabel metal1 2384 4562 2496 4578 0 _1235_.gnd
rlabel metal1 2384 4322 2496 4338 0 _1235_.vdd
rlabel metal2 2393 4493 2407 4507 0 _1235_.A
rlabel metal2 2413 4473 2427 4487 0 _1235_.B
rlabel metal2 2453 4453 2467 4467 0 _1235_.Y
rlabel metal1 2264 4562 2396 4578 0 _1195_.gnd
rlabel metal1 2264 4322 2396 4338 0 _1195_.vdd
rlabel metal2 2373 4473 2387 4487 0 _1195_.A
rlabel metal2 2353 4453 2367 4467 0 _1195_.B
rlabel metal2 2293 4473 2307 4487 0 _1195_.C
rlabel metal2 2333 4473 2347 4487 0 _1195_.Y
rlabel metal2 2313 4453 2327 4467 0 _1195_.D
rlabel metal1 2484 4562 2596 4578 0 _1236_.gnd
rlabel metal1 2484 4322 2596 4338 0 _1236_.vdd
rlabel metal2 2493 4453 2507 4467 0 _1236_.A
rlabel metal2 2513 4493 2527 4507 0 _1236_.B
rlabel metal2 2533 4453 2547 4467 0 _1236_.C
rlabel metal2 2553 4473 2567 4487 0 _1236_.Y
rlabel metal1 2584 4562 2716 4578 0 _1237_.gnd
rlabel metal1 2584 4322 2716 4338 0 _1237_.vdd
rlabel metal2 2693 4473 2707 4487 0 _1237_.A
rlabel metal2 2673 4453 2687 4467 0 _1237_.B
rlabel metal2 2613 4473 2627 4487 0 _1237_.C
rlabel metal2 2633 4453 2647 4467 0 _1237_.D
rlabel metal2 2653 4473 2667 4487 0 _1237_.Y
rlabel metal1 2704 4562 2956 4578 0 _1555_.gnd
rlabel metal1 2704 4322 2956 4338 0 _1555_.vdd
rlabel metal2 2793 4473 2807 4487 0 _1555_.D
rlabel metal2 2833 4473 2847 4487 0 _1555_.CLK
rlabel metal2 2913 4473 2927 4487 0 _1555_.Q
rlabel metal1 3184 4562 3296 4578 0 _1419_.gnd
rlabel metal1 3184 4322 3296 4338 0 _1419_.vdd
rlabel metal2 3273 4473 3287 4487 0 _1419_.A
rlabel metal2 3253 4453 3267 4467 0 _1419_.B
rlabel metal2 3213 4453 3227 4467 0 _1419_.C
rlabel metal2 3233 4473 3247 4487 0 _1419_.Y
rlabel metal1 3004 4562 3116 4578 0 _1418_.gnd
rlabel metal1 3004 4322 3116 4338 0 _1418_.vdd
rlabel metal2 3093 4473 3107 4487 0 _1418_.A
rlabel metal2 3073 4453 3087 4467 0 _1418_.B
rlabel metal2 3033 4453 3047 4467 0 _1418_.C
rlabel metal2 3053 4473 3067 4487 0 _1418_.Y
rlabel metal1 3104 4562 3196 4578 0 _1409_.gnd
rlabel metal1 3104 4322 3196 4338 0 _1409_.vdd
rlabel metal2 3133 4473 3147 4487 0 _1409_.B
rlabel metal2 3173 4473 3187 4487 0 _1409_.A
rlabel metal2 3153 4493 3167 4507 0 _1409_.Y
rlabel metal1 2944 4562 3016 4578 0 _1196_.gnd
rlabel metal1 2944 4322 3016 4338 0 _1196_.vdd
rlabel metal2 2993 4493 3007 4507 0 _1196_.A
rlabel metal2 2973 4453 2987 4467 0 _1196_.Y
rlabel metal1 3424 4562 3676 4578 0 _1539_.gnd
rlabel metal1 3424 4322 3676 4338 0 _1539_.vdd
rlabel metal2 3573 4473 3587 4487 0 _1539_.D
rlabel metal2 3533 4473 3547 4487 0 _1539_.CLK
rlabel metal2 3453 4473 3467 4487 0 _1539_.Q
rlabel metal1 3284 4562 3376 4578 0 _1410_.gnd
rlabel metal1 3284 4322 3376 4338 0 _1410_.vdd
rlabel metal2 3313 4473 3327 4487 0 _1410_.B
rlabel metal2 3353 4473 3367 4487 0 _1410_.A
rlabel metal2 3333 4493 3347 4507 0 _1410_.Y
rlabel metal1 3364 4562 3436 4578 0 _830_.gnd
rlabel metal1 3364 4322 3436 4338 0 _830_.vdd
rlabel metal2 3413 4493 3427 4507 0 _830_.A
rlabel metal2 3393 4453 3407 4467 0 _830_.Y
rlabel metal1 3664 4562 3776 4578 0 _832_.gnd
rlabel metal1 3664 4322 3776 4338 0 _832_.vdd
rlabel metal2 3673 4473 3687 4487 0 _832_.A
rlabel metal2 3693 4453 3707 4467 0 _832_.B
rlabel metal2 3733 4453 3747 4467 0 _832_.C
rlabel metal2 3713 4473 3727 4487 0 _832_.Y
rlabel metal1 3844 4562 4056 4578 0 CLKBUF1_insert10.gnd
rlabel metal1 3844 4322 4056 4338 0 CLKBUF1_insert10.vdd
rlabel metal2 4013 4453 4027 4467 0 CLKBUF1_insert10.A
rlabel metal2 3873 4453 3887 4467 0 CLKBUF1_insert10.Y
rlabel metal1 3764 4562 3856 4578 0 _831_.gnd
rlabel metal1 3764 4322 3856 4338 0 _831_.vdd
rlabel metal2 3773 4433 3787 4447 0 _831_.A
rlabel metal2 3813 4433 3827 4447 0 _831_.B
rlabel metal2 3793 4453 3807 4467 0 _831_.Y
rlabel metal1 4044 4562 4136 4578 0 _1601_.gnd
rlabel metal1 4044 4322 4136 4338 0 _1601_.vdd
rlabel metal2 4113 4473 4127 4487 0 _1601_.A
rlabel metal2 4073 4473 4087 4487 0 _1601_.Y
rlabel metal1 4264 4562 4376 4578 0 _838_.gnd
rlabel metal1 4264 4322 4376 4338 0 _838_.vdd
rlabel metal2 4273 4473 4287 4487 0 _838_.A
rlabel metal2 4293 4453 4307 4467 0 _838_.B
rlabel metal2 4333 4453 4347 4467 0 _838_.C
rlabel metal2 4313 4473 4327 4487 0 _838_.Y
rlabel metal1 4124 4562 4216 4578 0 _837_.gnd
rlabel metal1 4124 4322 4216 4338 0 _837_.vdd
rlabel metal2 4133 4433 4147 4447 0 _837_.A
rlabel metal2 4173 4433 4187 4447 0 _837_.B
rlabel metal2 4153 4453 4167 4467 0 _837_.Y
rlabel metal1 4204 4562 4276 4578 0 _836_.gnd
rlabel metal1 4204 4322 4276 4338 0 _836_.vdd
rlabel metal2 4213 4493 4227 4507 0 _836_.A
rlabel metal2 4233 4453 4247 4467 0 _836_.Y
rlabel metal1 4364 4562 4616 4578 0 _1541_.gnd
rlabel metal1 4364 4322 4616 4338 0 _1541_.vdd
rlabel metal2 4513 4473 4527 4487 0 _1541_.D
rlabel metal2 4473 4473 4487 4487 0 _1541_.CLK
rlabel metal2 4393 4473 4407 4487 0 _1541_.Q
rlabel metal1 4604 4562 4696 4578 0 _1609_.gnd
rlabel metal1 4604 4322 4696 4338 0 _1609_.vdd
rlabel metal2 4613 4473 4627 4487 0 _1609_.A
rlabel metal2 4653 4473 4667 4487 0 _1609_.Y
rlabel metal1 4684 4562 4776 4578 0 _1487_.gnd
rlabel metal1 4684 4322 4776 4338 0 _1487_.vdd
rlabel metal2 4693 4433 4707 4447 0 _1487_.A
rlabel metal2 4733 4433 4747 4447 0 _1487_.B
rlabel metal2 4713 4453 4727 4467 0 _1487_.Y
<< end >>
