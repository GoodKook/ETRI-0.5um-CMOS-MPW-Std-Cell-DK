magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 162 162
<< diffusion >>
rect 5 5 101 101
<< metal1 >>
rect 4 4 102 102
<< end >>
