magic
tech scmos
magscale 1 60
timestamp 1709340318
<< checkpaint >>
rect 6840 51320 10620 51360
rect -1210 51300 10620 51320
rect -1210 49320 11340 51300
rect -1210 49303 11710 49320
rect -2607 -3200 11710 49303
rect -2607 -3217 133 -3200
<< nwell >>
rect 310 42200 8410 45520
rect 310 22600 8410 38200
<< psubstratepdiff >>
rect 310 46800 8410 50120
rect 310 0 8410 15600
<< nsubstratendiff >>
rect 310 42200 8410 45520
rect 310 22600 8410 38200
<< metal1 >>
rect 310 46800 8410 50120
rect 310 42200 8410 45520
rect 310 22600 8410 38200
rect 310 0 8410 15600
<< metal2 >>
rect 310 46800 8410 50120
rect 310 42200 8410 45520
rect 310 22600 8410 38200
rect 310 0 8410 15600
<< metal3 >>
rect 310 46800 8410 50120
rect 310 42200 8410 45520
rect 310 22600 8410 38200
rect 310 0 8410 15600
use IOFILLER10  IOFILLER10_0
timestamp 1692859860
transform 1 0 70 0 1 0
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_1
timestamp 1692859860
transform 1 0 6650 0 1 0
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_2
timestamp 1692859860
transform 1 0 1710 0 1 0
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_3
timestamp 1692859860
transform 1 0 3350 0 1 0
box -70 0 2070 50120
use IOFILLER10  IOFILLER10_4
timestamp 1692859860
transform 1 0 5010 0 1 0
box -70 0 2070 50120
<< end >>
